.title 1-layer Power Grid for b04.points
* resistance segment model:
.subckt Rseg 1 3
R1 1 2 0.583
L1 2 3 0.003n
C1 1 0 0.25e-12
C2 3 0 0.25e-12
.ends
* the horizontal resistors:
X1 n_40280_40040 n_40660_40040 Rseg
X2 n_40660_40040 n_41420_40040 Rseg
X3 n_41420_40040 n_41800_40040 Rseg
X4 n_41800_40040 n_42180_40040 Rseg
X5 n_42180_40040 n_42940_40040 Rseg
X6 n_42940_40040 n_43320_40040 Rseg
X7 n_43320_40040 n_43700_40040 Rseg
X8 n_43700_40040 n_44080_40040 Rseg
X9 n_44080_40040 n_44460_40040 Rseg
X10 n_44460_40040 n_44840_40040 Rseg
X11 n_44840_40040 n_45220_40040 Rseg
X12 n_45220_40040 n_45600_40040 Rseg
X13 n_45600_40040 n_46360_40040 Rseg
X14 n_46360_40040 n_46740_40040 Rseg
X15 n_46740_40040 n_47120_40040 Rseg
X16 n_47120_40040 n_47500_40040 Rseg
X17 n_47500_40040 n_47880_40040 Rseg
X18 n_47880_40040 n_48260_40040 Rseg
X19 n_48260_40040 n_48640_40040 Rseg
X20 n_48640_40040 n_49020_40040 Rseg
X21 n_49020_40040 n_49400_40040 Rseg
X22 n_49400_40040 n_49780_40040 Rseg
X23 n_49780_40040 n_50160_40040 Rseg
X24 n_50160_40040 n_50540_40040 Rseg
X25 n_50540_40040 n_50920_40040 Rseg
X26 n_50920_40040 n_51300_40040 Rseg
X27 n_51300_40040 n_51680_40040 Rseg
X28 n_51680_40040 n_52060_40040 Rseg
X29 n_52060_40040 n_52440_40040 Rseg
X30 n_52440_40040 n_52820_40040 Rseg
X31 n_52820_40040 n_53200_40040 Rseg
X32 n_53200_40040 n_53580_40040 Rseg
X33 n_53580_40040 n_53960_40040 Rseg
X34 n_53960_40040 n_54340_40040 Rseg
X35 n_54340_40040 n_54720_40040 Rseg
X36 n_54720_40040 n_55100_40040 Rseg
X37 n_55100_40040 n_55480_40040 Rseg
X38 n_55480_40040 n_55860_40040 Rseg
X39 n_55860_40040 n_56240_40040 Rseg
X40 n_56240_40040 n_56620_40040 Rseg
X41 n_56620_40040 n_57000_40040 Rseg
X42 n_57000_40040 n_57380_40040 Rseg
X43 n_57380_40040 n_57760_40040 Rseg
X44 n_57760_40040 n_58140_40040 Rseg
X45 n_58140_40040 n_58520_40040 Rseg
X46 n_58520_40040 n_58900_40040 Rseg
X47 n_58900_40040 n_59280_40040 Rseg
X48 n_59280_40040 n_59660_40040 Rseg
X49 n_59660_40040 n_60040_40040 Rseg
X50 n_60040_40040 n_60420_40040 Rseg
X51 n_60420_40040 n_60800_40040 Rseg
X52 n_60800_40040 n_61180_40040 Rseg
X53 n_61180_40040 n_61560_40040 Rseg
X54 n_61560_40040 n_61940_40040 Rseg
X55 n_61940_40040 n_62320_40040 Rseg
X56 n_62320_40040 n_63080_40040 Rseg
X57 n_63080_40040 n_63460_40040 Rseg
X58 n_63460_40040 n_63840_40040 Rseg
X59 n_63840_40040 n_64220_40040 Rseg
X60 n_64220_40040 n_64600_40040 Rseg
X61 n_64600_40040 n_64980_40040 Rseg
X62 n_64980_40040 n_65360_40040 Rseg
X63 n_65360_40040 n_65740_40040 Rseg
X64 n_65740_40040 n_66120_40040 Rseg
X65 n_66120_40040 n_66880_40040 Rseg
X66 n_66880_40040 n_67260_40040 Rseg
X67 n_67260_40040 n_68020_40040 Rseg
X68 n_68020_40040 n_68400_40040 Rseg
X69 n_68400_40040 n_68780_40040 Rseg
X70 n_68780_40040 n_69160_40040 Rseg
X71 n_69160_40040 n_69920_40040 Rseg
X72 n_69920_40040 n_70300_40040 Rseg
X73 n_70300_40040 n_71060_40040 Rseg
X74 n_71060_40040 n_71820_40040 Rseg
X75 n_71820_40040 n_72200_40040 Rseg
X76 n_72200_40040 n_72960_40040 Rseg
X77 n_72960_40040 n_73340_40040 Rseg
X78 n_73340_40040 n_73720_40040 Rseg
X79 n_73720_40040 n_74100_40040 Rseg
X80 n_74100_40040 n_74860_40040 Rseg
X81 n_74860_40040 n_75240_40040 Rseg
X82 n_75240_40040 n_76000_40040 Rseg
X83 n_76000_40040 n_76380_40040 Rseg
X84 n_76380_40040 n_76760_40040 Rseg
X85 n_76760_40040 n_77140_40040 Rseg
X86 n_77140_40040 n_77520_40040 Rseg
X87 n_77520_40040 n_77900_40040 Rseg
X88 n_77900_40040 n_78280_40040 Rseg
X89 n_78280_40040 n_78660_40040 Rseg
X90 n_78660_40040 n_79040_40040 Rseg
X91 n_79040_40040 n_80180_40040 Rseg
X92 n_80180_40040 n_80560_40040 Rseg
X93 n_80560_40040 n_80940_40040 Rseg
X94 n_80940_40040 n_81700_40040 Rseg
X95 n_81700_40040 n_82080_40040 Rseg
X96 n_82080_40040 n_83220_40040 Rseg
X97 n_83220_40040 n_83600_40040 Rseg
X98 n_83600_40040 n_84740_40040 Rseg
X99 n_84740_40040 n_85120_40040 Rseg
X100 n_85120_40040 n_85500_40040 Rseg
X101 n_85500_40040 n_85880_40040 Rseg
X102 n_85880_40040 n_86260_40040 Rseg
X103 n_86260_40040 n_87020_40040 Rseg
X104 n_87020_40040 n_87400_40040 Rseg
X105 n_87400_40040 n_87780_40040 Rseg
X106 n_87780_40040 n_88160_40040 Rseg
X107 n_88160_40040 n_88540_40040 Rseg
X108 n_88540_40040 n_88920_40040 Rseg
X109 n_88920_40040 n_89300_40040 Rseg
X110 n_89300_40040 n_90060_40040 Rseg
X111 n_90060_40040 n_90440_40040 Rseg
X112 n_90440_40040 n_90820_40040 Rseg
X113 n_90820_40040 n_91200_40040 Rseg
X114 n_91200_40040 n_91580_40040 Rseg
X115 n_91580_40040 n_91960_40040 Rseg
X116 n_91960_40040 n_92340_40040 Rseg
X117 n_92340_40040 n_92720_40040 Rseg
X118 n_92720_40040 n_93100_40040 Rseg
X119 n_93100_40040 n_93480_40040 Rseg
X120 n_40280_42840 n_40660_42840 Rseg
X121 n_40660_42840 n_41420_42840 Rseg
X122 n_41420_42840 n_41800_42840 Rseg
X123 n_41800_42840 n_42180_42840 Rseg
X124 n_42180_42840 n_42940_42840 Rseg
X125 n_42940_42840 n_43320_42840 Rseg
X126 n_43320_42840 n_43700_42840 Rseg
X127 n_43700_42840 n_44080_42840 Rseg
X128 n_44080_42840 n_44460_42840 Rseg
X129 n_44460_42840 n_44840_42840 Rseg
X130 n_44840_42840 n_45220_42840 Rseg
X131 n_45220_42840 n_45600_42840 Rseg
X132 n_45600_42840 n_46360_42840 Rseg
X133 n_46360_42840 n_46740_42840 Rseg
X134 n_46740_42840 n_47120_42840 Rseg
X135 n_47120_42840 n_47500_42840 Rseg
X136 n_47500_42840 n_47880_42840 Rseg
X137 n_47880_42840 n_48260_42840 Rseg
X138 n_48260_42840 n_48640_42840 Rseg
X139 n_48640_42840 n_49020_42840 Rseg
X140 n_49020_42840 n_49400_42840 Rseg
X141 n_49400_42840 n_49780_42840 Rseg
X142 n_49780_42840 n_50160_42840 Rseg
X143 n_50160_42840 n_50540_42840 Rseg
X144 n_50540_42840 n_50920_42840 Rseg
X145 n_50920_42840 n_51300_42840 Rseg
X146 n_51300_42840 n_51680_42840 Rseg
X147 n_51680_42840 n_52060_42840 Rseg
X148 n_52060_42840 n_52440_42840 Rseg
X149 n_52440_42840 n_52820_42840 Rseg
X150 n_52820_42840 n_53200_42840 Rseg
X151 n_53200_42840 n_53580_42840 Rseg
X152 n_53580_42840 n_53960_42840 Rseg
X153 n_53960_42840 n_54340_42840 Rseg
X154 n_54340_42840 n_54720_42840 Rseg
X155 n_54720_42840 n_55100_42840 Rseg
X156 n_55100_42840 n_55480_42840 Rseg
X157 n_55480_42840 n_55860_42840 Rseg
X158 n_55860_42840 n_56240_42840 Rseg
X159 n_56240_42840 n_56620_42840 Rseg
X160 n_56620_42840 n_57000_42840 Rseg
X161 n_57000_42840 n_57380_42840 Rseg
X162 n_57380_42840 n_57760_42840 Rseg
X163 n_57760_42840 n_58140_42840 Rseg
X164 n_58140_42840 n_58520_42840 Rseg
X165 n_58520_42840 n_58900_42840 Rseg
X166 n_58900_42840 n_59280_42840 Rseg
X167 n_59280_42840 n_59660_42840 Rseg
X168 n_59660_42840 n_60040_42840 Rseg
X169 n_60040_42840 n_60420_42840 Rseg
X170 n_60420_42840 n_60800_42840 Rseg
X171 n_60800_42840 n_61180_42840 Rseg
X172 n_61180_42840 n_61560_42840 Rseg
X173 n_61560_42840 n_61940_42840 Rseg
X174 n_61940_42840 n_62320_42840 Rseg
X175 n_62320_42840 n_63080_42840 Rseg
X176 n_63080_42840 n_63460_42840 Rseg
X177 n_63460_42840 n_63840_42840 Rseg
X178 n_63840_42840 n_64220_42840 Rseg
X179 n_64220_42840 n_64600_42840 Rseg
X180 n_64600_42840 n_64980_42840 Rseg
X181 n_64980_42840 n_65360_42840 Rseg
X182 n_65360_42840 n_65740_42840 Rseg
X183 n_65740_42840 n_66120_42840 Rseg
X184 n_66120_42840 n_66880_42840 Rseg
X185 n_66880_42840 n_67260_42840 Rseg
X186 n_67260_42840 n_68020_42840 Rseg
X187 n_68020_42840 n_68400_42840 Rseg
X188 n_68400_42840 n_68780_42840 Rseg
X189 n_68780_42840 n_69160_42840 Rseg
X190 n_69160_42840 n_69920_42840 Rseg
X191 n_69920_42840 n_70300_42840 Rseg
X192 n_70300_42840 n_71060_42840 Rseg
X193 n_71060_42840 n_71820_42840 Rseg
X194 n_71820_42840 n_72200_42840 Rseg
X195 n_72200_42840 n_72960_42840 Rseg
X196 n_72960_42840 n_73340_42840 Rseg
X197 n_73340_42840 n_73720_42840 Rseg
X198 n_73720_42840 n_74100_42840 Rseg
X199 n_74100_42840 n_74860_42840 Rseg
X200 n_74860_42840 n_75240_42840 Rseg
X201 n_75240_42840 n_76000_42840 Rseg
X202 n_76000_42840 n_76380_42840 Rseg
X203 n_76380_42840 n_76760_42840 Rseg
X204 n_76760_42840 n_77140_42840 Rseg
X205 n_77140_42840 n_77520_42840 Rseg
X206 n_77520_42840 n_77900_42840 Rseg
X207 n_77900_42840 n_78280_42840 Rseg
X208 n_78280_42840 n_78660_42840 Rseg
X209 n_78660_42840 n_79040_42840 Rseg
X210 n_79040_42840 n_80180_42840 Rseg
X211 n_80180_42840 n_80560_42840 Rseg
X212 n_80560_42840 n_80940_42840 Rseg
X213 n_80940_42840 n_81700_42840 Rseg
X214 n_81700_42840 n_82080_42840 Rseg
X215 n_82080_42840 n_83220_42840 Rseg
X216 n_83220_42840 n_83600_42840 Rseg
X217 n_83600_42840 n_84740_42840 Rseg
X218 n_84740_42840 n_85120_42840 Rseg
X219 n_85120_42840 n_85500_42840 Rseg
X220 n_85500_42840 n_85880_42840 Rseg
X221 n_85880_42840 n_86260_42840 Rseg
X222 n_86260_42840 n_87020_42840 Rseg
X223 n_87020_42840 n_87400_42840 Rseg
X224 n_87400_42840 n_87780_42840 Rseg
X225 n_87780_42840 n_88160_42840 Rseg
X226 n_88160_42840 n_88540_42840 Rseg
X227 n_88540_42840 n_88920_42840 Rseg
X228 n_88920_42840 n_89300_42840 Rseg
X229 n_89300_42840 n_90060_42840 Rseg
X230 n_90060_42840 n_90440_42840 Rseg
X231 n_90440_42840 n_90820_42840 Rseg
X232 n_90820_42840 n_91200_42840 Rseg
X233 n_91200_42840 n_91580_42840 Rseg
X234 n_91580_42840 n_91960_42840 Rseg
X235 n_91960_42840 n_92340_42840 Rseg
X236 n_92340_42840 n_92720_42840 Rseg
X237 n_92720_42840 n_93100_42840 Rseg
X238 n_93100_42840 n_93480_42840 Rseg
X239 n_40280_45640 n_40660_45640 Rseg
X240 n_40660_45640 n_41420_45640 Rseg
X241 n_41420_45640 n_41800_45640 Rseg
X242 n_41800_45640 n_42180_45640 Rseg
X243 n_42180_45640 n_42940_45640 Rseg
X244 n_42940_45640 n_43320_45640 Rseg
X245 n_43320_45640 n_43700_45640 Rseg
X246 n_43700_45640 n_44080_45640 Rseg
X247 n_44080_45640 n_44460_45640 Rseg
X248 n_44460_45640 n_44840_45640 Rseg
X249 n_44840_45640 n_45220_45640 Rseg
X250 n_45220_45640 n_45600_45640 Rseg
X251 n_45600_45640 n_46360_45640 Rseg
X252 n_46360_45640 n_46740_45640 Rseg
X253 n_46740_45640 n_47120_45640 Rseg
X254 n_47120_45640 n_47500_45640 Rseg
X255 n_47500_45640 n_47880_45640 Rseg
X256 n_47880_45640 n_48260_45640 Rseg
X257 n_48260_45640 n_48640_45640 Rseg
X258 n_48640_45640 n_49020_45640 Rseg
X259 n_49020_45640 n_49400_45640 Rseg
X260 n_49400_45640 n_49780_45640 Rseg
X261 n_49780_45640 n_50160_45640 Rseg
X262 n_50160_45640 n_50540_45640 Rseg
X263 n_50540_45640 n_50920_45640 Rseg
X264 n_50920_45640 n_51300_45640 Rseg
X265 n_51300_45640 n_51680_45640 Rseg
X266 n_51680_45640 n_52060_45640 Rseg
X267 n_52060_45640 n_52440_45640 Rseg
X268 n_52440_45640 n_52820_45640 Rseg
X269 n_52820_45640 n_53200_45640 Rseg
X270 n_53200_45640 n_53580_45640 Rseg
X271 n_53580_45640 n_53960_45640 Rseg
X272 n_53960_45640 n_54340_45640 Rseg
X273 n_54340_45640 n_54720_45640 Rseg
X274 n_54720_45640 n_55100_45640 Rseg
X275 n_55100_45640 n_55480_45640 Rseg
X276 n_55480_45640 n_55860_45640 Rseg
X277 n_55860_45640 n_56240_45640 Rseg
X278 n_56240_45640 n_56620_45640 Rseg
X279 n_56620_45640 n_57000_45640 Rseg
X280 n_57000_45640 n_57380_45640 Rseg
X281 n_57380_45640 n_57760_45640 Rseg
X282 n_57760_45640 n_58140_45640 Rseg
X283 n_58140_45640 n_58520_45640 Rseg
X284 n_58520_45640 n_58900_45640 Rseg
X285 n_58900_45640 n_59280_45640 Rseg
X286 n_59280_45640 n_59660_45640 Rseg
X287 n_59660_45640 n_60040_45640 Rseg
X288 n_60040_45640 n_60420_45640 Rseg
X289 n_60420_45640 n_60800_45640 Rseg
X290 n_60800_45640 n_61180_45640 Rseg
X291 n_61180_45640 n_61560_45640 Rseg
X292 n_61560_45640 n_61940_45640 Rseg
X293 n_61940_45640 n_62320_45640 Rseg
X294 n_62320_45640 n_63080_45640 Rseg
X295 n_63080_45640 n_63460_45640 Rseg
X296 n_63460_45640 n_63840_45640 Rseg
X297 n_63840_45640 n_64220_45640 Rseg
X298 n_64220_45640 n_64600_45640 Rseg
X299 n_64600_45640 n_64980_45640 Rseg
X300 n_64980_45640 n_65360_45640 Rseg
X301 n_65360_45640 n_65740_45640 Rseg
X302 n_65740_45640 n_66120_45640 Rseg
X303 n_66120_45640 n_66880_45640 Rseg
X304 n_66880_45640 n_67260_45640 Rseg
X305 n_67260_45640 n_68020_45640 Rseg
X306 n_68020_45640 n_68400_45640 Rseg
X307 n_68400_45640 n_68780_45640 Rseg
X308 n_68780_45640 n_69160_45640 Rseg
X309 n_69160_45640 n_69920_45640 Rseg
X310 n_69920_45640 n_70300_45640 Rseg
X311 n_70300_45640 n_71060_45640 Rseg
X312 n_71060_45640 n_71820_45640 Rseg
X313 n_71820_45640 n_72200_45640 Rseg
X314 n_72200_45640 n_72960_45640 Rseg
X315 n_72960_45640 n_73340_45640 Rseg
X316 n_73340_45640 n_73720_45640 Rseg
X317 n_73720_45640 n_74100_45640 Rseg
X318 n_74100_45640 n_74860_45640 Rseg
X319 n_74860_45640 n_75240_45640 Rseg
X320 n_75240_45640 n_76000_45640 Rseg
X321 n_76000_45640 n_76380_45640 Rseg
X322 n_76380_45640 n_76760_45640 Rseg
X323 n_76760_45640 n_77140_45640 Rseg
X324 n_77140_45640 n_77520_45640 Rseg
X325 n_77520_45640 n_77900_45640 Rseg
X326 n_77900_45640 n_78280_45640 Rseg
X327 n_78280_45640 n_78660_45640 Rseg
X328 n_78660_45640 n_79040_45640 Rseg
X329 n_79040_45640 n_80180_45640 Rseg
X330 n_80180_45640 n_80560_45640 Rseg
X331 n_80560_45640 n_80940_45640 Rseg
X332 n_80940_45640 n_81700_45640 Rseg
X333 n_81700_45640 n_82080_45640 Rseg
X334 n_82080_45640 n_83220_45640 Rseg
X335 n_83220_45640 n_83600_45640 Rseg
X336 n_83600_45640 n_84740_45640 Rseg
X337 n_84740_45640 n_85120_45640 Rseg
X338 n_85120_45640 n_85500_45640 Rseg
X339 n_85500_45640 n_85880_45640 Rseg
X340 n_85880_45640 n_86260_45640 Rseg
X341 n_86260_45640 n_87020_45640 Rseg
X342 n_87020_45640 n_87400_45640 Rseg
X343 n_87400_45640 n_87780_45640 Rseg
X344 n_87780_45640 n_88160_45640 Rseg
X345 n_88160_45640 n_88540_45640 Rseg
X346 n_88540_45640 n_88920_45640 Rseg
X347 n_88920_45640 n_89300_45640 Rseg
X348 n_89300_45640 n_90060_45640 Rseg
X349 n_90060_45640 n_90440_45640 Rseg
X350 n_90440_45640 n_90820_45640 Rseg
X351 n_90820_45640 n_91200_45640 Rseg
X352 n_91200_45640 n_91580_45640 Rseg
X353 n_91580_45640 n_91960_45640 Rseg
X354 n_91960_45640 n_92340_45640 Rseg
X355 n_92340_45640 n_92720_45640 Rseg
X356 n_92720_45640 n_93100_45640 Rseg
X357 n_93100_45640 n_93480_45640 Rseg
X358 n_40280_48440 n_40660_48440 Rseg
X359 n_40660_48440 n_41420_48440 Rseg
X360 n_41420_48440 n_41800_48440 Rseg
X361 n_41800_48440 n_42180_48440 Rseg
X362 n_42180_48440 n_42940_48440 Rseg
X363 n_42940_48440 n_43320_48440 Rseg
X364 n_43320_48440 n_43700_48440 Rseg
X365 n_43700_48440 n_44080_48440 Rseg
X366 n_44080_48440 n_44460_48440 Rseg
X367 n_44460_48440 n_44840_48440 Rseg
X368 n_44840_48440 n_45220_48440 Rseg
X369 n_45220_48440 n_45600_48440 Rseg
X370 n_45600_48440 n_46360_48440 Rseg
X371 n_46360_48440 n_46740_48440 Rseg
X372 n_46740_48440 n_47120_48440 Rseg
X373 n_47120_48440 n_47500_48440 Rseg
X374 n_47500_48440 n_47880_48440 Rseg
X375 n_47880_48440 n_48260_48440 Rseg
X376 n_48260_48440 n_48640_48440 Rseg
X377 n_48640_48440 n_49020_48440 Rseg
X378 n_49020_48440 n_49400_48440 Rseg
X379 n_49400_48440 n_49780_48440 Rseg
X380 n_49780_48440 n_50160_48440 Rseg
X381 n_50160_48440 n_50540_48440 Rseg
X382 n_50540_48440 n_50920_48440 Rseg
X383 n_50920_48440 n_51300_48440 Rseg
X384 n_51300_48440 n_51680_48440 Rseg
X385 n_51680_48440 n_52060_48440 Rseg
X386 n_52060_48440 n_52440_48440 Rseg
X387 n_52440_48440 n_52820_48440 Rseg
X388 n_52820_48440 n_53200_48440 Rseg
X389 n_53200_48440 n_53580_48440 Rseg
X390 n_53580_48440 n_53960_48440 Rseg
X391 n_53960_48440 n_54340_48440 Rseg
X392 n_54340_48440 n_54720_48440 Rseg
X393 n_54720_48440 n_55100_48440 Rseg
X394 n_55100_48440 n_55480_48440 Rseg
X395 n_55480_48440 n_55860_48440 Rseg
X396 n_55860_48440 n_56240_48440 Rseg
X397 n_56240_48440 n_56620_48440 Rseg
X398 n_56620_48440 n_57000_48440 Rseg
X399 n_57000_48440 n_57380_48440 Rseg
X400 n_57380_48440 n_57760_48440 Rseg
X401 n_57760_48440 n_58140_48440 Rseg
X402 n_58140_48440 n_58520_48440 Rseg
X403 n_58520_48440 n_58900_48440 Rseg
X404 n_58900_48440 n_59280_48440 Rseg
X405 n_59280_48440 n_59660_48440 Rseg
X406 n_59660_48440 n_60040_48440 Rseg
X407 n_60040_48440 n_60420_48440 Rseg
X408 n_60420_48440 n_60800_48440 Rseg
X409 n_60800_48440 n_61180_48440 Rseg
X410 n_61180_48440 n_61560_48440 Rseg
X411 n_61560_48440 n_61940_48440 Rseg
X412 n_61940_48440 n_62320_48440 Rseg
X413 n_62320_48440 n_63080_48440 Rseg
X414 n_63080_48440 n_63460_48440 Rseg
X415 n_63460_48440 n_63840_48440 Rseg
X416 n_63840_48440 n_64220_48440 Rseg
X417 n_64220_48440 n_64600_48440 Rseg
X418 n_64600_48440 n_64980_48440 Rseg
X419 n_64980_48440 n_65360_48440 Rseg
X420 n_65360_48440 n_65740_48440 Rseg
X421 n_65740_48440 n_66120_48440 Rseg
X422 n_66120_48440 n_66880_48440 Rseg
X423 n_66880_48440 n_67260_48440 Rseg
X424 n_67260_48440 n_68020_48440 Rseg
X425 n_68020_48440 n_68400_48440 Rseg
X426 n_68400_48440 n_68780_48440 Rseg
X427 n_68780_48440 n_69160_48440 Rseg
X428 n_69160_48440 n_69920_48440 Rseg
X429 n_69920_48440 n_70300_48440 Rseg
X430 n_70300_48440 n_71060_48440 Rseg
X431 n_71060_48440 n_71820_48440 Rseg
X432 n_71820_48440 n_72200_48440 Rseg
X433 n_72200_48440 n_72960_48440 Rseg
X434 n_72960_48440 n_73340_48440 Rseg
X435 n_73340_48440 n_73720_48440 Rseg
X436 n_73720_48440 n_74100_48440 Rseg
X437 n_74100_48440 n_74860_48440 Rseg
X438 n_74860_48440 n_75240_48440 Rseg
X439 n_75240_48440 n_76000_48440 Rseg
X440 n_76000_48440 n_76380_48440 Rseg
X441 n_76380_48440 n_76760_48440 Rseg
X442 n_76760_48440 n_77140_48440 Rseg
X443 n_77140_48440 n_77520_48440 Rseg
X444 n_77520_48440 n_77900_48440 Rseg
X445 n_77900_48440 n_78280_48440 Rseg
X446 n_78280_48440 n_78660_48440 Rseg
X447 n_78660_48440 n_79040_48440 Rseg
X448 n_79040_48440 n_80180_48440 Rseg
X449 n_80180_48440 n_80560_48440 Rseg
X450 n_80560_48440 n_80940_48440 Rseg
X451 n_80940_48440 n_81700_48440 Rseg
X452 n_81700_48440 n_82080_48440 Rseg
X453 n_82080_48440 n_83220_48440 Rseg
X454 n_83220_48440 n_83600_48440 Rseg
X455 n_83600_48440 n_84740_48440 Rseg
X456 n_84740_48440 n_85120_48440 Rseg
X457 n_85120_48440 n_85500_48440 Rseg
X458 n_85500_48440 n_85880_48440 Rseg
X459 n_85880_48440 n_86260_48440 Rseg
X460 n_86260_48440 n_87020_48440 Rseg
X461 n_87020_48440 n_87400_48440 Rseg
X462 n_87400_48440 n_87780_48440 Rseg
X463 n_87780_48440 n_88160_48440 Rseg
X464 n_88160_48440 n_88540_48440 Rseg
X465 n_88540_48440 n_88920_48440 Rseg
X466 n_88920_48440 n_89300_48440 Rseg
X467 n_89300_48440 n_90060_48440 Rseg
X468 n_90060_48440 n_90440_48440 Rseg
X469 n_90440_48440 n_90820_48440 Rseg
X470 n_90820_48440 n_91200_48440 Rseg
X471 n_91200_48440 n_91580_48440 Rseg
X472 n_91580_48440 n_91960_48440 Rseg
X473 n_91960_48440 n_92340_48440 Rseg
X474 n_92340_48440 n_92720_48440 Rseg
X475 n_92720_48440 n_93100_48440 Rseg
X476 n_93100_48440 n_93480_48440 Rseg
X477 n_40280_51240 n_40660_51240 Rseg
X478 n_40660_51240 n_41420_51240 Rseg
X479 n_41420_51240 n_41800_51240 Rseg
X480 n_41800_51240 n_42180_51240 Rseg
X481 n_42180_51240 n_42940_51240 Rseg
X482 n_42940_51240 n_43320_51240 Rseg
X483 n_43320_51240 n_43700_51240 Rseg
X484 n_43700_51240 n_44080_51240 Rseg
X485 n_44080_51240 n_44460_51240 Rseg
X486 n_44460_51240 n_44840_51240 Rseg
X487 n_44840_51240 n_45220_51240 Rseg
X488 n_45220_51240 n_45600_51240 Rseg
X489 n_45600_51240 n_46360_51240 Rseg
X490 n_46360_51240 n_46740_51240 Rseg
X491 n_46740_51240 n_47120_51240 Rseg
X492 n_47120_51240 n_47500_51240 Rseg
X493 n_47500_51240 n_47880_51240 Rseg
X494 n_47880_51240 n_48260_51240 Rseg
X495 n_48260_51240 n_48640_51240 Rseg
X496 n_48640_51240 n_49020_51240 Rseg
X497 n_49020_51240 n_49400_51240 Rseg
X498 n_49400_51240 n_49780_51240 Rseg
X499 n_49780_51240 n_50160_51240 Rseg
X500 n_50160_51240 n_50540_51240 Rseg
X501 n_50540_51240 n_50920_51240 Rseg
X502 n_50920_51240 n_51300_51240 Rseg
X503 n_51300_51240 n_51680_51240 Rseg
X504 n_51680_51240 n_52060_51240 Rseg
X505 n_52060_51240 n_52440_51240 Rseg
X506 n_52440_51240 n_52820_51240 Rseg
X507 n_52820_51240 n_53200_51240 Rseg
X508 n_53200_51240 n_53580_51240 Rseg
X509 n_53580_51240 n_53960_51240 Rseg
X510 n_53960_51240 n_54340_51240 Rseg
X511 n_54340_51240 n_54720_51240 Rseg
X512 n_54720_51240 n_55100_51240 Rseg
X513 n_55100_51240 n_55480_51240 Rseg
X514 n_55480_51240 n_55860_51240 Rseg
X515 n_55860_51240 n_56240_51240 Rseg
X516 n_56240_51240 n_56620_51240 Rseg
X517 n_56620_51240 n_57000_51240 Rseg
X518 n_57000_51240 n_57380_51240 Rseg
X519 n_57380_51240 n_57760_51240 Rseg
X520 n_57760_51240 n_58140_51240 Rseg
X521 n_58140_51240 n_58520_51240 Rseg
X522 n_58520_51240 n_58900_51240 Rseg
X523 n_58900_51240 n_59280_51240 Rseg
X524 n_59280_51240 n_59660_51240 Rseg
X525 n_59660_51240 n_60040_51240 Rseg
X526 n_60040_51240 n_60420_51240 Rseg
X527 n_60420_51240 n_60800_51240 Rseg
X528 n_60800_51240 n_61180_51240 Rseg
X529 n_61180_51240 n_61560_51240 Rseg
X530 n_61560_51240 n_61940_51240 Rseg
X531 n_61940_51240 n_62320_51240 Rseg
X532 n_62320_51240 n_63080_51240 Rseg
X533 n_63080_51240 n_63460_51240 Rseg
X534 n_63460_51240 n_63840_51240 Rseg
X535 n_63840_51240 n_64220_51240 Rseg
X536 n_64220_51240 n_64600_51240 Rseg
X537 n_64600_51240 n_64980_51240 Rseg
X538 n_64980_51240 n_65360_51240 Rseg
X539 n_65360_51240 n_65740_51240 Rseg
X540 n_65740_51240 n_66120_51240 Rseg
X541 n_66120_51240 n_66880_51240 Rseg
X542 n_66880_51240 n_67260_51240 Rseg
X543 n_67260_51240 n_68020_51240 Rseg
X544 n_68020_51240 n_68400_51240 Rseg
X545 n_68400_51240 n_68780_51240 Rseg
X546 n_68780_51240 n_69160_51240 Rseg
X547 n_69160_51240 n_69920_51240 Rseg
X548 n_69920_51240 n_70300_51240 Rseg
X549 n_70300_51240 n_71060_51240 Rseg
X550 n_71060_51240 n_71820_51240 Rseg
X551 n_71820_51240 n_72200_51240 Rseg
X552 n_72200_51240 n_72960_51240 Rseg
X553 n_72960_51240 n_73340_51240 Rseg
X554 n_73340_51240 n_73720_51240 Rseg
X555 n_73720_51240 n_74100_51240 Rseg
X556 n_74100_51240 n_74860_51240 Rseg
X557 n_74860_51240 n_75240_51240 Rseg
X558 n_75240_51240 n_76000_51240 Rseg
X559 n_76000_51240 n_76380_51240 Rseg
X560 n_76380_51240 n_76760_51240 Rseg
X561 n_76760_51240 n_77140_51240 Rseg
X562 n_77140_51240 n_77520_51240 Rseg
X563 n_77520_51240 n_77900_51240 Rseg
X564 n_77900_51240 n_78280_51240 Rseg
X565 n_78280_51240 n_78660_51240 Rseg
X566 n_78660_51240 n_79040_51240 Rseg
X567 n_79040_51240 n_80180_51240 Rseg
X568 n_80180_51240 n_80560_51240 Rseg
X569 n_80560_51240 n_80940_51240 Rseg
X570 n_80940_51240 n_81700_51240 Rseg
X571 n_81700_51240 n_82080_51240 Rseg
X572 n_82080_51240 n_83220_51240 Rseg
X573 n_83220_51240 n_83600_51240 Rseg
X574 n_83600_51240 n_84740_51240 Rseg
X575 n_84740_51240 n_85120_51240 Rseg
X576 n_85120_51240 n_85500_51240 Rseg
X577 n_85500_51240 n_85880_51240 Rseg
X578 n_85880_51240 n_86260_51240 Rseg
X579 n_86260_51240 n_87020_51240 Rseg
X580 n_87020_51240 n_87400_51240 Rseg
X581 n_87400_51240 n_87780_51240 Rseg
X582 n_87780_51240 n_88160_51240 Rseg
X583 n_88160_51240 n_88540_51240 Rseg
X584 n_88540_51240 n_88920_51240 Rseg
X585 n_88920_51240 n_89300_51240 Rseg
X586 n_89300_51240 n_90060_51240 Rseg
X587 n_90060_51240 n_90440_51240 Rseg
X588 n_90440_51240 n_90820_51240 Rseg
X589 n_90820_51240 n_91200_51240 Rseg
X590 n_91200_51240 n_91580_51240 Rseg
X591 n_91580_51240 n_91960_51240 Rseg
X592 n_91960_51240 n_92340_51240 Rseg
X593 n_92340_51240 n_92720_51240 Rseg
X594 n_92720_51240 n_93100_51240 Rseg
X595 n_93100_51240 n_93480_51240 Rseg
X596 n_40280_54040 n_40660_54040 Rseg
X597 n_40660_54040 n_41420_54040 Rseg
X598 n_41420_54040 n_41800_54040 Rseg
X599 n_41800_54040 n_42180_54040 Rseg
X600 n_42180_54040 n_42940_54040 Rseg
X601 n_42940_54040 n_43320_54040 Rseg
X602 n_43320_54040 n_43700_54040 Rseg
X603 n_43700_54040 n_44080_54040 Rseg
X604 n_44080_54040 n_44460_54040 Rseg
X605 n_44460_54040 n_44840_54040 Rseg
X606 n_44840_54040 n_45220_54040 Rseg
X607 n_45220_54040 n_45600_54040 Rseg
X608 n_45600_54040 n_46360_54040 Rseg
X609 n_46360_54040 n_46740_54040 Rseg
X610 n_46740_54040 n_47120_54040 Rseg
X611 n_47120_54040 n_47500_54040 Rseg
X612 n_47500_54040 n_47880_54040 Rseg
X613 n_47880_54040 n_48260_54040 Rseg
X614 n_48260_54040 n_48640_54040 Rseg
X615 n_48640_54040 n_49020_54040 Rseg
X616 n_49020_54040 n_49400_54040 Rseg
X617 n_49400_54040 n_49780_54040 Rseg
X618 n_49780_54040 n_50160_54040 Rseg
X619 n_50160_54040 n_50540_54040 Rseg
X620 n_50540_54040 n_50920_54040 Rseg
X621 n_50920_54040 n_51300_54040 Rseg
X622 n_51300_54040 n_51680_54040 Rseg
X623 n_51680_54040 n_52060_54040 Rseg
X624 n_52060_54040 n_52440_54040 Rseg
X625 n_52440_54040 n_52820_54040 Rseg
X626 n_52820_54040 n_53200_54040 Rseg
X627 n_53200_54040 n_53580_54040 Rseg
X628 n_53580_54040 n_53960_54040 Rseg
X629 n_53960_54040 n_54340_54040 Rseg
X630 n_54340_54040 n_54720_54040 Rseg
X631 n_54720_54040 n_55100_54040 Rseg
X632 n_55100_54040 n_55480_54040 Rseg
X633 n_55480_54040 n_55860_54040 Rseg
X634 n_55860_54040 n_56240_54040 Rseg
X635 n_56240_54040 n_56620_54040 Rseg
X636 n_56620_54040 n_57000_54040 Rseg
X637 n_57000_54040 n_57380_54040 Rseg
X638 n_57380_54040 n_57760_54040 Rseg
X639 n_57760_54040 n_58140_54040 Rseg
X640 n_58140_54040 n_58520_54040 Rseg
X641 n_58520_54040 n_58900_54040 Rseg
X642 n_58900_54040 n_59280_54040 Rseg
X643 n_59280_54040 n_59660_54040 Rseg
X644 n_59660_54040 n_60040_54040 Rseg
X645 n_60040_54040 n_60420_54040 Rseg
X646 n_60420_54040 n_60800_54040 Rseg
X647 n_60800_54040 n_61180_54040 Rseg
X648 n_61180_54040 n_61560_54040 Rseg
X649 n_61560_54040 n_61940_54040 Rseg
X650 n_61940_54040 n_62320_54040 Rseg
X651 n_62320_54040 n_63080_54040 Rseg
X652 n_63080_54040 n_63460_54040 Rseg
X653 n_63460_54040 n_63840_54040 Rseg
X654 n_63840_54040 n_64220_54040 Rseg
X655 n_64220_54040 n_64600_54040 Rseg
X656 n_64600_54040 n_64980_54040 Rseg
X657 n_64980_54040 n_65360_54040 Rseg
X658 n_65360_54040 n_65740_54040 Rseg
X659 n_65740_54040 n_66120_54040 Rseg
X660 n_66120_54040 n_66880_54040 Rseg
X661 n_66880_54040 n_67260_54040 Rseg
X662 n_67260_54040 n_68020_54040 Rseg
X663 n_68020_54040 n_68400_54040 Rseg
X664 n_68400_54040 n_68780_54040 Rseg
X665 n_68780_54040 n_69160_54040 Rseg
X666 n_69160_54040 n_69920_54040 Rseg
X667 n_69920_54040 n_70300_54040 Rseg
X668 n_70300_54040 n_71060_54040 Rseg
X669 n_71060_54040 n_71820_54040 Rseg
X670 n_71820_54040 n_72200_54040 Rseg
X671 n_72200_54040 n_72960_54040 Rseg
X672 n_72960_54040 n_73340_54040 Rseg
X673 n_73340_54040 n_73720_54040 Rseg
X674 n_73720_54040 n_74100_54040 Rseg
X675 n_74100_54040 n_74860_54040 Rseg
X676 n_74860_54040 n_75240_54040 Rseg
X677 n_75240_54040 n_76000_54040 Rseg
X678 n_76000_54040 n_76380_54040 Rseg
X679 n_76380_54040 n_76760_54040 Rseg
X680 n_76760_54040 n_77140_54040 Rseg
X681 n_77140_54040 n_77520_54040 Rseg
X682 n_77520_54040 n_77900_54040 Rseg
X683 n_77900_54040 n_78280_54040 Rseg
X684 n_78280_54040 n_78660_54040 Rseg
X685 n_78660_54040 n_79040_54040 Rseg
X686 n_79040_54040 n_80180_54040 Rseg
X687 n_80180_54040 n_80560_54040 Rseg
X688 n_80560_54040 n_80940_54040 Rseg
X689 n_80940_54040 n_81700_54040 Rseg
X690 n_81700_54040 n_82080_54040 Rseg
X691 n_82080_54040 n_83220_54040 Rseg
X692 n_83220_54040 n_83600_54040 Rseg
X693 n_83600_54040 n_84740_54040 Rseg
X694 n_84740_54040 n_85120_54040 Rseg
X695 n_85120_54040 n_85500_54040 Rseg
X696 n_85500_54040 n_85880_54040 Rseg
X697 n_85880_54040 n_86260_54040 Rseg
X698 n_86260_54040 n_87020_54040 Rseg
X699 n_87020_54040 n_87400_54040 Rseg
X700 n_87400_54040 n_87780_54040 Rseg
X701 n_87780_54040 n_88160_54040 Rseg
X702 n_88160_54040 n_88540_54040 Rseg
X703 n_88540_54040 n_88920_54040 Rseg
X704 n_88920_54040 n_89300_54040 Rseg
X705 n_89300_54040 n_90060_54040 Rseg
X706 n_90060_54040 n_90440_54040 Rseg
X707 n_90440_54040 n_90820_54040 Rseg
X708 n_90820_54040 n_91200_54040 Rseg
X709 n_91200_54040 n_91580_54040 Rseg
X710 n_91580_54040 n_91960_54040 Rseg
X711 n_91960_54040 n_92340_54040 Rseg
X712 n_92340_54040 n_92720_54040 Rseg
X713 n_92720_54040 n_93100_54040 Rseg
X714 n_93100_54040 n_93480_54040 Rseg
X715 n_40280_56840 n_40660_56840 Rseg
X716 n_40660_56840 n_41420_56840 Rseg
X717 n_41420_56840 n_41800_56840 Rseg
X718 n_41800_56840 n_42180_56840 Rseg
X719 n_42180_56840 n_42940_56840 Rseg
X720 n_42940_56840 n_43320_56840 Rseg
X721 n_43320_56840 n_43700_56840 Rseg
X722 n_43700_56840 n_44080_56840 Rseg
X723 n_44080_56840 n_44460_56840 Rseg
X724 n_44460_56840 n_44840_56840 Rseg
X725 n_44840_56840 n_45220_56840 Rseg
X726 n_45220_56840 n_45600_56840 Rseg
X727 n_45600_56840 n_46360_56840 Rseg
X728 n_46360_56840 n_46740_56840 Rseg
X729 n_46740_56840 n_47120_56840 Rseg
X730 n_47120_56840 n_47500_56840 Rseg
X731 n_47500_56840 n_47880_56840 Rseg
X732 n_47880_56840 n_48260_56840 Rseg
X733 n_48260_56840 n_48640_56840 Rseg
X734 n_48640_56840 n_49020_56840 Rseg
X735 n_49020_56840 n_49400_56840 Rseg
X736 n_49400_56840 n_49780_56840 Rseg
X737 n_49780_56840 n_50160_56840 Rseg
X738 n_50160_56840 n_50540_56840 Rseg
X739 n_50540_56840 n_50920_56840 Rseg
X740 n_50920_56840 n_51300_56840 Rseg
X741 n_51300_56840 n_51680_56840 Rseg
X742 n_51680_56840 n_52060_56840 Rseg
X743 n_52060_56840 n_52440_56840 Rseg
X744 n_52440_56840 n_52820_56840 Rseg
X745 n_52820_56840 n_53200_56840 Rseg
X746 n_53200_56840 n_53580_56840 Rseg
X747 n_53580_56840 n_53960_56840 Rseg
X748 n_53960_56840 n_54340_56840 Rseg
X749 n_54340_56840 n_54720_56840 Rseg
X750 n_54720_56840 n_55100_56840 Rseg
X751 n_55100_56840 n_55480_56840 Rseg
X752 n_55480_56840 n_55860_56840 Rseg
X753 n_55860_56840 n_56240_56840 Rseg
X754 n_56240_56840 n_56620_56840 Rseg
X755 n_56620_56840 n_57000_56840 Rseg
X756 n_57000_56840 n_57380_56840 Rseg
X757 n_57380_56840 n_57760_56840 Rseg
X758 n_57760_56840 n_58140_56840 Rseg
X759 n_58140_56840 n_58520_56840 Rseg
X760 n_58520_56840 n_58900_56840 Rseg
X761 n_58900_56840 n_59280_56840 Rseg
X762 n_59280_56840 n_59660_56840 Rseg
X763 n_59660_56840 n_60040_56840 Rseg
X764 n_60040_56840 n_60420_56840 Rseg
X765 n_60420_56840 n_60800_56840 Rseg
X766 n_60800_56840 n_61180_56840 Rseg
X767 n_61180_56840 n_61560_56840 Rseg
X768 n_61560_56840 n_61940_56840 Rseg
X769 n_61940_56840 n_62320_56840 Rseg
X770 n_62320_56840 n_63080_56840 Rseg
X771 n_63080_56840 n_63460_56840 Rseg
X772 n_63460_56840 n_63840_56840 Rseg
X773 n_63840_56840 n_64220_56840 Rseg
X774 n_64220_56840 n_64600_56840 Rseg
X775 n_64600_56840 n_64980_56840 Rseg
X776 n_64980_56840 n_65360_56840 Rseg
X777 n_65360_56840 n_65740_56840 Rseg
X778 n_65740_56840 n_66120_56840 Rseg
X779 n_66120_56840 n_66880_56840 Rseg
X780 n_66880_56840 n_67260_56840 Rseg
X781 n_67260_56840 n_68020_56840 Rseg
X782 n_68020_56840 n_68400_56840 Rseg
X783 n_68400_56840 n_68780_56840 Rseg
X784 n_68780_56840 n_69160_56840 Rseg
X785 n_69160_56840 n_69920_56840 Rseg
X786 n_69920_56840 n_70300_56840 Rseg
X787 n_70300_56840 n_71060_56840 Rseg
X788 n_71060_56840 n_71820_56840 Rseg
X789 n_71820_56840 n_72200_56840 Rseg
X790 n_72200_56840 n_72960_56840 Rseg
X791 n_72960_56840 n_73340_56840 Rseg
X792 n_73340_56840 n_73720_56840 Rseg
X793 n_73720_56840 n_74100_56840 Rseg
X794 n_74100_56840 n_74860_56840 Rseg
X795 n_74860_56840 n_75240_56840 Rseg
X796 n_75240_56840 n_76000_56840 Rseg
X797 n_76000_56840 n_76380_56840 Rseg
X798 n_76380_56840 n_76760_56840 Rseg
X799 n_76760_56840 n_77140_56840 Rseg
X800 n_77140_56840 n_77520_56840 Rseg
X801 n_77520_56840 n_77900_56840 Rseg
X802 n_77900_56840 n_78280_56840 Rseg
X803 n_78280_56840 n_78660_56840 Rseg
X804 n_78660_56840 n_79040_56840 Rseg
X805 n_79040_56840 n_80180_56840 Rseg
X806 n_80180_56840 n_80560_56840 Rseg
X807 n_80560_56840 n_80940_56840 Rseg
X808 n_80940_56840 n_81700_56840 Rseg
X809 n_81700_56840 n_82080_56840 Rseg
X810 n_82080_56840 n_83220_56840 Rseg
X811 n_83220_56840 n_83600_56840 Rseg
X812 n_83600_56840 n_84740_56840 Rseg
X813 n_84740_56840 n_85120_56840 Rseg
X814 n_85120_56840 n_85500_56840 Rseg
X815 n_85500_56840 n_85880_56840 Rseg
X816 n_85880_56840 n_86260_56840 Rseg
X817 n_86260_56840 n_87020_56840 Rseg
X818 n_87020_56840 n_87400_56840 Rseg
X819 n_87400_56840 n_87780_56840 Rseg
X820 n_87780_56840 n_88160_56840 Rseg
X821 n_88160_56840 n_88540_56840 Rseg
X822 n_88540_56840 n_88920_56840 Rseg
X823 n_88920_56840 n_89300_56840 Rseg
X824 n_89300_56840 n_90060_56840 Rseg
X825 n_90060_56840 n_90440_56840 Rseg
X826 n_90440_56840 n_90820_56840 Rseg
X827 n_90820_56840 n_91200_56840 Rseg
X828 n_91200_56840 n_91580_56840 Rseg
X829 n_91580_56840 n_91960_56840 Rseg
X830 n_91960_56840 n_92340_56840 Rseg
X831 n_92340_56840 n_92720_56840 Rseg
X832 n_92720_56840 n_93100_56840 Rseg
X833 n_93100_56840 n_93480_56840 Rseg
X834 n_40280_59640 n_40660_59640 Rseg
X835 n_40660_59640 n_41420_59640 Rseg
X836 n_41420_59640 n_41800_59640 Rseg
X837 n_41800_59640 n_42180_59640 Rseg
X838 n_42180_59640 n_42940_59640 Rseg
X839 n_42940_59640 n_43320_59640 Rseg
X840 n_43320_59640 n_43700_59640 Rseg
X841 n_43700_59640 n_44080_59640 Rseg
X842 n_44080_59640 n_44460_59640 Rseg
X843 n_44460_59640 n_44840_59640 Rseg
X844 n_44840_59640 n_45220_59640 Rseg
X845 n_45220_59640 n_45600_59640 Rseg
X846 n_45600_59640 n_46360_59640 Rseg
X847 n_46360_59640 n_46740_59640 Rseg
X848 n_46740_59640 n_47120_59640 Rseg
X849 n_47120_59640 n_47500_59640 Rseg
X850 n_47500_59640 n_47880_59640 Rseg
X851 n_47880_59640 n_48260_59640 Rseg
X852 n_48260_59640 n_48640_59640 Rseg
X853 n_48640_59640 n_49020_59640 Rseg
X854 n_49020_59640 n_49400_59640 Rseg
X855 n_49400_59640 n_49780_59640 Rseg
X856 n_49780_59640 n_50160_59640 Rseg
X857 n_50160_59640 n_50540_59640 Rseg
X858 n_50540_59640 n_50920_59640 Rseg
X859 n_50920_59640 n_51300_59640 Rseg
X860 n_51300_59640 n_51680_59640 Rseg
X861 n_51680_59640 n_52060_59640 Rseg
X862 n_52060_59640 n_52440_59640 Rseg
X863 n_52440_59640 n_52820_59640 Rseg
X864 n_52820_59640 n_53200_59640 Rseg
X865 n_53200_59640 n_53580_59640 Rseg
X866 n_53580_59640 n_53960_59640 Rseg
X867 n_53960_59640 n_54340_59640 Rseg
X868 n_54340_59640 n_54720_59640 Rseg
X869 n_54720_59640 n_55100_59640 Rseg
X870 n_55100_59640 n_55480_59640 Rseg
X871 n_55480_59640 n_55860_59640 Rseg
X872 n_55860_59640 n_56240_59640 Rseg
X873 n_56240_59640 n_56620_59640 Rseg
X874 n_56620_59640 n_57000_59640 Rseg
X875 n_57000_59640 n_57380_59640 Rseg
X876 n_57380_59640 n_57760_59640 Rseg
X877 n_57760_59640 n_58140_59640 Rseg
X878 n_58140_59640 n_58520_59640 Rseg
X879 n_58520_59640 n_58900_59640 Rseg
X880 n_58900_59640 n_59280_59640 Rseg
X881 n_59280_59640 n_59660_59640 Rseg
X882 n_59660_59640 n_60040_59640 Rseg
X883 n_60040_59640 n_60420_59640 Rseg
X884 n_60420_59640 n_60800_59640 Rseg
X885 n_60800_59640 n_61180_59640 Rseg
X886 n_61180_59640 n_61560_59640 Rseg
X887 n_61560_59640 n_61940_59640 Rseg
X888 n_61940_59640 n_62320_59640 Rseg
X889 n_62320_59640 n_63080_59640 Rseg
X890 n_63080_59640 n_63460_59640 Rseg
X891 n_63460_59640 n_63840_59640 Rseg
X892 n_63840_59640 n_64220_59640 Rseg
X893 n_64220_59640 n_64600_59640 Rseg
X894 n_64600_59640 n_64980_59640 Rseg
X895 n_64980_59640 n_65360_59640 Rseg
X896 n_65360_59640 n_65740_59640 Rseg
X897 n_65740_59640 n_66120_59640 Rseg
X898 n_66120_59640 n_66880_59640 Rseg
X899 n_66880_59640 n_67260_59640 Rseg
X900 n_67260_59640 n_68020_59640 Rseg
X901 n_68020_59640 n_68400_59640 Rseg
X902 n_68400_59640 n_68780_59640 Rseg
X903 n_68780_59640 n_69160_59640 Rseg
X904 n_69160_59640 n_69920_59640 Rseg
X905 n_69920_59640 n_70300_59640 Rseg
X906 n_70300_59640 n_71060_59640 Rseg
X907 n_71060_59640 n_71820_59640 Rseg
X908 n_71820_59640 n_72200_59640 Rseg
X909 n_72200_59640 n_72960_59640 Rseg
X910 n_72960_59640 n_73340_59640 Rseg
X911 n_73340_59640 n_73720_59640 Rseg
X912 n_73720_59640 n_74100_59640 Rseg
X913 n_74100_59640 n_74860_59640 Rseg
X914 n_74860_59640 n_75240_59640 Rseg
X915 n_75240_59640 n_76000_59640 Rseg
X916 n_76000_59640 n_76380_59640 Rseg
X917 n_76380_59640 n_76760_59640 Rseg
X918 n_76760_59640 n_77140_59640 Rseg
X919 n_77140_59640 n_77520_59640 Rseg
X920 n_77520_59640 n_77900_59640 Rseg
X921 n_77900_59640 n_78280_59640 Rseg
X922 n_78280_59640 n_78660_59640 Rseg
X923 n_78660_59640 n_79040_59640 Rseg
X924 n_79040_59640 n_80180_59640 Rseg
X925 n_80180_59640 n_80560_59640 Rseg
X926 n_80560_59640 n_80940_59640 Rseg
X927 n_80940_59640 n_81700_59640 Rseg
X928 n_81700_59640 n_82080_59640 Rseg
X929 n_82080_59640 n_83220_59640 Rseg
X930 n_83220_59640 n_83600_59640 Rseg
X931 n_83600_59640 n_84740_59640 Rseg
X932 n_84740_59640 n_85120_59640 Rseg
X933 n_85120_59640 n_85500_59640 Rseg
X934 n_85500_59640 n_85880_59640 Rseg
X935 n_85880_59640 n_86260_59640 Rseg
X936 n_86260_59640 n_87020_59640 Rseg
X937 n_87020_59640 n_87400_59640 Rseg
X938 n_87400_59640 n_87780_59640 Rseg
X939 n_87780_59640 n_88160_59640 Rseg
X940 n_88160_59640 n_88540_59640 Rseg
X941 n_88540_59640 n_88920_59640 Rseg
X942 n_88920_59640 n_89300_59640 Rseg
X943 n_89300_59640 n_90060_59640 Rseg
X944 n_90060_59640 n_90440_59640 Rseg
X945 n_90440_59640 n_90820_59640 Rseg
X946 n_90820_59640 n_91200_59640 Rseg
X947 n_91200_59640 n_91580_59640 Rseg
X948 n_91580_59640 n_91960_59640 Rseg
X949 n_91960_59640 n_92340_59640 Rseg
X950 n_92340_59640 n_92720_59640 Rseg
X951 n_92720_59640 n_93100_59640 Rseg
X952 n_93100_59640 n_93480_59640 Rseg
X953 n_40280_62440 n_40660_62440 Rseg
X954 n_40660_62440 n_41420_62440 Rseg
X955 n_41420_62440 n_41800_62440 Rseg
X956 n_41800_62440 n_42180_62440 Rseg
X957 n_42180_62440 n_42940_62440 Rseg
X958 n_42940_62440 n_43320_62440 Rseg
X959 n_43320_62440 n_43700_62440 Rseg
X960 n_43700_62440 n_44080_62440 Rseg
X961 n_44080_62440 n_44460_62440 Rseg
X962 n_44460_62440 n_44840_62440 Rseg
X963 n_44840_62440 n_45220_62440 Rseg
X964 n_45220_62440 n_45600_62440 Rseg
X965 n_45600_62440 n_46360_62440 Rseg
X966 n_46360_62440 n_46740_62440 Rseg
X967 n_46740_62440 n_47120_62440 Rseg
X968 n_47120_62440 n_47500_62440 Rseg
X969 n_47500_62440 n_47880_62440 Rseg
X970 n_47880_62440 n_48260_62440 Rseg
X971 n_48260_62440 n_48640_62440 Rseg
X972 n_48640_62440 n_49020_62440 Rseg
X973 n_49020_62440 n_49400_62440 Rseg
X974 n_49400_62440 n_49780_62440 Rseg
X975 n_49780_62440 n_50160_62440 Rseg
X976 n_50160_62440 n_50540_62440 Rseg
X977 n_50540_62440 n_50920_62440 Rseg
X978 n_50920_62440 n_51300_62440 Rseg
X979 n_51300_62440 n_51680_62440 Rseg
X980 n_51680_62440 n_52060_62440 Rseg
X981 n_52060_62440 n_52440_62440 Rseg
X982 n_52440_62440 n_52820_62440 Rseg
X983 n_52820_62440 n_53200_62440 Rseg
X984 n_53200_62440 n_53580_62440 Rseg
X985 n_53580_62440 n_53960_62440 Rseg
X986 n_53960_62440 n_54340_62440 Rseg
X987 n_54340_62440 n_54720_62440 Rseg
X988 n_54720_62440 n_55100_62440 Rseg
X989 n_55100_62440 n_55480_62440 Rseg
X990 n_55480_62440 n_55860_62440 Rseg
X991 n_55860_62440 n_56240_62440 Rseg
X992 n_56240_62440 n_56620_62440 Rseg
X993 n_56620_62440 n_57000_62440 Rseg
X994 n_57000_62440 n_57380_62440 Rseg
X995 n_57380_62440 n_57760_62440 Rseg
X996 n_57760_62440 n_58140_62440 Rseg
X997 n_58140_62440 n_58520_62440 Rseg
X998 n_58520_62440 n_58900_62440 Rseg
X999 n_58900_62440 n_59280_62440 Rseg
X1000 n_59280_62440 n_59660_62440 Rseg
X1001 n_59660_62440 n_60040_62440 Rseg
X1002 n_60040_62440 n_60420_62440 Rseg
X1003 n_60420_62440 n_60800_62440 Rseg
X1004 n_60800_62440 n_61180_62440 Rseg
X1005 n_61180_62440 n_61560_62440 Rseg
X1006 n_61560_62440 n_61940_62440 Rseg
X1007 n_61940_62440 n_62320_62440 Rseg
X1008 n_62320_62440 n_63080_62440 Rseg
X1009 n_63080_62440 n_63460_62440 Rseg
X1010 n_63460_62440 n_63840_62440 Rseg
X1011 n_63840_62440 n_64220_62440 Rseg
X1012 n_64220_62440 n_64600_62440 Rseg
X1013 n_64600_62440 n_64980_62440 Rseg
X1014 n_64980_62440 n_65360_62440 Rseg
X1015 n_65360_62440 n_65740_62440 Rseg
X1016 n_65740_62440 n_66120_62440 Rseg
X1017 n_66120_62440 n_66880_62440 Rseg
X1018 n_66880_62440 n_67260_62440 Rseg
X1019 n_67260_62440 n_68020_62440 Rseg
X1020 n_68020_62440 n_68400_62440 Rseg
X1021 n_68400_62440 n_68780_62440 Rseg
X1022 n_68780_62440 n_69160_62440 Rseg
X1023 n_69160_62440 n_69920_62440 Rseg
X1024 n_69920_62440 n_70300_62440 Rseg
X1025 n_70300_62440 n_71060_62440 Rseg
X1026 n_71060_62440 n_71820_62440 Rseg
X1027 n_71820_62440 n_72200_62440 Rseg
X1028 n_72200_62440 n_72960_62440 Rseg
X1029 n_72960_62440 n_73340_62440 Rseg
X1030 n_73340_62440 n_73720_62440 Rseg
X1031 n_73720_62440 n_74100_62440 Rseg
X1032 n_74100_62440 n_74860_62440 Rseg
X1033 n_74860_62440 n_75240_62440 Rseg
X1034 n_75240_62440 n_76000_62440 Rseg
X1035 n_76000_62440 n_76380_62440 Rseg
X1036 n_76380_62440 n_76760_62440 Rseg
X1037 n_76760_62440 n_77140_62440 Rseg
X1038 n_77140_62440 n_77520_62440 Rseg
X1039 n_77520_62440 n_77900_62440 Rseg
X1040 n_77900_62440 n_78280_62440 Rseg
X1041 n_78280_62440 n_78660_62440 Rseg
X1042 n_78660_62440 n_79040_62440 Rseg
X1043 n_79040_62440 n_80180_62440 Rseg
X1044 n_80180_62440 n_80560_62440 Rseg
X1045 n_80560_62440 n_80940_62440 Rseg
X1046 n_80940_62440 n_81700_62440 Rseg
X1047 n_81700_62440 n_82080_62440 Rseg
X1048 n_82080_62440 n_83220_62440 Rseg
X1049 n_83220_62440 n_83600_62440 Rseg
X1050 n_83600_62440 n_84740_62440 Rseg
X1051 n_84740_62440 n_85120_62440 Rseg
X1052 n_85120_62440 n_85500_62440 Rseg
X1053 n_85500_62440 n_85880_62440 Rseg
X1054 n_85880_62440 n_86260_62440 Rseg
X1055 n_86260_62440 n_87020_62440 Rseg
X1056 n_87020_62440 n_87400_62440 Rseg
X1057 n_87400_62440 n_87780_62440 Rseg
X1058 n_87780_62440 n_88160_62440 Rseg
X1059 n_88160_62440 n_88540_62440 Rseg
X1060 n_88540_62440 n_88920_62440 Rseg
X1061 n_88920_62440 n_89300_62440 Rseg
X1062 n_89300_62440 n_90060_62440 Rseg
X1063 n_90060_62440 n_90440_62440 Rseg
X1064 n_90440_62440 n_90820_62440 Rseg
X1065 n_90820_62440 n_91200_62440 Rseg
X1066 n_91200_62440 n_91580_62440 Rseg
X1067 n_91580_62440 n_91960_62440 Rseg
X1068 n_91960_62440 n_92340_62440 Rseg
X1069 n_92340_62440 n_92720_62440 Rseg
X1070 n_92720_62440 n_93100_62440 Rseg
X1071 n_93100_62440 n_93480_62440 Rseg
X1072 n_40280_65240 n_40660_65240 Rseg
X1073 n_40660_65240 n_41420_65240 Rseg
X1074 n_41420_65240 n_41800_65240 Rseg
X1075 n_41800_65240 n_42180_65240 Rseg
X1076 n_42180_65240 n_42940_65240 Rseg
X1077 n_42940_65240 n_43320_65240 Rseg
X1078 n_43320_65240 n_43700_65240 Rseg
X1079 n_43700_65240 n_44080_65240 Rseg
X1080 n_44080_65240 n_44460_65240 Rseg
X1081 n_44460_65240 n_44840_65240 Rseg
X1082 n_44840_65240 n_45220_65240 Rseg
X1083 n_45220_65240 n_45600_65240 Rseg
X1084 n_45600_65240 n_46360_65240 Rseg
X1085 n_46360_65240 n_46740_65240 Rseg
X1086 n_46740_65240 n_47120_65240 Rseg
X1087 n_47120_65240 n_47500_65240 Rseg
X1088 n_47500_65240 n_47880_65240 Rseg
X1089 n_47880_65240 n_48260_65240 Rseg
X1090 n_48260_65240 n_48640_65240 Rseg
X1091 n_48640_65240 n_49020_65240 Rseg
X1092 n_49020_65240 n_49400_65240 Rseg
X1093 n_49400_65240 n_49780_65240 Rseg
X1094 n_49780_65240 n_50160_65240 Rseg
X1095 n_50160_65240 n_50540_65240 Rseg
X1096 n_50540_65240 n_50920_65240 Rseg
X1097 n_50920_65240 n_51300_65240 Rseg
X1098 n_51300_65240 n_51680_65240 Rseg
X1099 n_51680_65240 n_52060_65240 Rseg
X1100 n_52060_65240 n_52440_65240 Rseg
X1101 n_52440_65240 n_52820_65240 Rseg
X1102 n_52820_65240 n_53200_65240 Rseg
X1103 n_53200_65240 n_53580_65240 Rseg
X1104 n_53580_65240 n_53960_65240 Rseg
X1105 n_53960_65240 n_54340_65240 Rseg
X1106 n_54340_65240 n_54720_65240 Rseg
X1107 n_54720_65240 n_55100_65240 Rseg
X1108 n_55100_65240 n_55480_65240 Rseg
X1109 n_55480_65240 n_55860_65240 Rseg
X1110 n_55860_65240 n_56240_65240 Rseg
X1111 n_56240_65240 n_56620_65240 Rseg
X1112 n_56620_65240 n_57000_65240 Rseg
X1113 n_57000_65240 n_57380_65240 Rseg
X1114 n_57380_65240 n_57760_65240 Rseg
X1115 n_57760_65240 n_58140_65240 Rseg
X1116 n_58140_65240 n_58520_65240 Rseg
X1117 n_58520_65240 n_58900_65240 Rseg
X1118 n_58900_65240 n_59280_65240 Rseg
X1119 n_59280_65240 n_59660_65240 Rseg
X1120 n_59660_65240 n_60040_65240 Rseg
X1121 n_60040_65240 n_60420_65240 Rseg
X1122 n_60420_65240 n_60800_65240 Rseg
X1123 n_60800_65240 n_61180_65240 Rseg
X1124 n_61180_65240 n_61560_65240 Rseg
X1125 n_61560_65240 n_61940_65240 Rseg
X1126 n_61940_65240 n_62320_65240 Rseg
X1127 n_62320_65240 n_63080_65240 Rseg
X1128 n_63080_65240 n_63460_65240 Rseg
X1129 n_63460_65240 n_63840_65240 Rseg
X1130 n_63840_65240 n_64220_65240 Rseg
X1131 n_64220_65240 n_64600_65240 Rseg
X1132 n_64600_65240 n_64980_65240 Rseg
X1133 n_64980_65240 n_65360_65240 Rseg
X1134 n_65360_65240 n_65740_65240 Rseg
X1135 n_65740_65240 n_66120_65240 Rseg
X1136 n_66120_65240 n_66880_65240 Rseg
X1137 n_66880_65240 n_67260_65240 Rseg
X1138 n_67260_65240 n_68020_65240 Rseg
X1139 n_68020_65240 n_68400_65240 Rseg
X1140 n_68400_65240 n_68780_65240 Rseg
X1141 n_68780_65240 n_69160_65240 Rseg
X1142 n_69160_65240 n_69920_65240 Rseg
X1143 n_69920_65240 n_70300_65240 Rseg
X1144 n_70300_65240 n_71060_65240 Rseg
X1145 n_71060_65240 n_71820_65240 Rseg
X1146 n_71820_65240 n_72200_65240 Rseg
X1147 n_72200_65240 n_72960_65240 Rseg
X1148 n_72960_65240 n_73340_65240 Rseg
X1149 n_73340_65240 n_73720_65240 Rseg
X1150 n_73720_65240 n_74100_65240 Rseg
X1151 n_74100_65240 n_74860_65240 Rseg
X1152 n_74860_65240 n_75240_65240 Rseg
X1153 n_75240_65240 n_76000_65240 Rseg
X1154 n_76000_65240 n_76380_65240 Rseg
X1155 n_76380_65240 n_76760_65240 Rseg
X1156 n_76760_65240 n_77140_65240 Rseg
X1157 n_77140_65240 n_77520_65240 Rseg
X1158 n_77520_65240 n_77900_65240 Rseg
X1159 n_77900_65240 n_78280_65240 Rseg
X1160 n_78280_65240 n_78660_65240 Rseg
X1161 n_78660_65240 n_79040_65240 Rseg
X1162 n_79040_65240 n_80180_65240 Rseg
X1163 n_80180_65240 n_80560_65240 Rseg
X1164 n_80560_65240 n_80940_65240 Rseg
X1165 n_80940_65240 n_81700_65240 Rseg
X1166 n_81700_65240 n_82080_65240 Rseg
X1167 n_82080_65240 n_83220_65240 Rseg
X1168 n_83220_65240 n_83600_65240 Rseg
X1169 n_83600_65240 n_84740_65240 Rseg
X1170 n_84740_65240 n_85120_65240 Rseg
X1171 n_85120_65240 n_85500_65240 Rseg
X1172 n_85500_65240 n_85880_65240 Rseg
X1173 n_85880_65240 n_86260_65240 Rseg
X1174 n_86260_65240 n_87020_65240 Rseg
X1175 n_87020_65240 n_87400_65240 Rseg
X1176 n_87400_65240 n_87780_65240 Rseg
X1177 n_87780_65240 n_88160_65240 Rseg
X1178 n_88160_65240 n_88540_65240 Rseg
X1179 n_88540_65240 n_88920_65240 Rseg
X1180 n_88920_65240 n_89300_65240 Rseg
X1181 n_89300_65240 n_90060_65240 Rseg
X1182 n_90060_65240 n_90440_65240 Rseg
X1183 n_90440_65240 n_90820_65240 Rseg
X1184 n_90820_65240 n_91200_65240 Rseg
X1185 n_91200_65240 n_91580_65240 Rseg
X1186 n_91580_65240 n_91960_65240 Rseg
X1187 n_91960_65240 n_92340_65240 Rseg
X1188 n_92340_65240 n_92720_65240 Rseg
X1189 n_92720_65240 n_93100_65240 Rseg
X1190 n_93100_65240 n_93480_65240 Rseg
X1191 n_40280_68040 n_40660_68040 Rseg
X1192 n_40660_68040 n_41420_68040 Rseg
X1193 n_41420_68040 n_41800_68040 Rseg
X1194 n_41800_68040 n_42180_68040 Rseg
X1195 n_42180_68040 n_42940_68040 Rseg
X1196 n_42940_68040 n_43320_68040 Rseg
X1197 n_43320_68040 n_43700_68040 Rseg
X1198 n_43700_68040 n_44080_68040 Rseg
X1199 n_44080_68040 n_44460_68040 Rseg
X1200 n_44460_68040 n_44840_68040 Rseg
X1201 n_44840_68040 n_45220_68040 Rseg
X1202 n_45220_68040 n_45600_68040 Rseg
X1203 n_45600_68040 n_46360_68040 Rseg
X1204 n_46360_68040 n_46740_68040 Rseg
X1205 n_46740_68040 n_47120_68040 Rseg
X1206 n_47120_68040 n_47500_68040 Rseg
X1207 n_47500_68040 n_47880_68040 Rseg
X1208 n_47880_68040 n_48260_68040 Rseg
X1209 n_48260_68040 n_48640_68040 Rseg
X1210 n_48640_68040 n_49020_68040 Rseg
X1211 n_49020_68040 n_49400_68040 Rseg
X1212 n_49400_68040 n_49780_68040 Rseg
X1213 n_49780_68040 n_50160_68040 Rseg
X1214 n_50160_68040 n_50540_68040 Rseg
X1215 n_50540_68040 n_50920_68040 Rseg
X1216 n_50920_68040 n_51300_68040 Rseg
X1217 n_51300_68040 n_51680_68040 Rseg
X1218 n_51680_68040 n_52060_68040 Rseg
X1219 n_52060_68040 n_52440_68040 Rseg
X1220 n_52440_68040 n_52820_68040 Rseg
X1221 n_52820_68040 n_53200_68040 Rseg
X1222 n_53200_68040 n_53580_68040 Rseg
X1223 n_53580_68040 n_53960_68040 Rseg
X1224 n_53960_68040 n_54340_68040 Rseg
X1225 n_54340_68040 n_54720_68040 Rseg
X1226 n_54720_68040 n_55100_68040 Rseg
X1227 n_55100_68040 n_55480_68040 Rseg
X1228 n_55480_68040 n_55860_68040 Rseg
X1229 n_55860_68040 n_56240_68040 Rseg
X1230 n_56240_68040 n_56620_68040 Rseg
X1231 n_56620_68040 n_57000_68040 Rseg
X1232 n_57000_68040 n_57380_68040 Rseg
X1233 n_57380_68040 n_57760_68040 Rseg
X1234 n_57760_68040 n_58140_68040 Rseg
X1235 n_58140_68040 n_58520_68040 Rseg
X1236 n_58520_68040 n_58900_68040 Rseg
X1237 n_58900_68040 n_59280_68040 Rseg
X1238 n_59280_68040 n_59660_68040 Rseg
X1239 n_59660_68040 n_60040_68040 Rseg
X1240 n_60040_68040 n_60420_68040 Rseg
X1241 n_60420_68040 n_60800_68040 Rseg
X1242 n_60800_68040 n_61180_68040 Rseg
X1243 n_61180_68040 n_61560_68040 Rseg
X1244 n_61560_68040 n_61940_68040 Rseg
X1245 n_61940_68040 n_62320_68040 Rseg
X1246 n_62320_68040 n_63080_68040 Rseg
X1247 n_63080_68040 n_63460_68040 Rseg
X1248 n_63460_68040 n_63840_68040 Rseg
X1249 n_63840_68040 n_64220_68040 Rseg
X1250 n_64220_68040 n_64600_68040 Rseg
X1251 n_64600_68040 n_64980_68040 Rseg
X1252 n_64980_68040 n_65360_68040 Rseg
X1253 n_65360_68040 n_65740_68040 Rseg
X1254 n_65740_68040 n_66120_68040 Rseg
X1255 n_66120_68040 n_66880_68040 Rseg
X1256 n_66880_68040 n_67260_68040 Rseg
X1257 n_67260_68040 n_68020_68040 Rseg
X1258 n_68020_68040 n_68400_68040 Rseg
X1259 n_68400_68040 n_68780_68040 Rseg
X1260 n_68780_68040 n_69160_68040 Rseg
X1261 n_69160_68040 n_69920_68040 Rseg
X1262 n_69920_68040 n_70300_68040 Rseg
X1263 n_70300_68040 n_71060_68040 Rseg
X1264 n_71060_68040 n_71820_68040 Rseg
X1265 n_71820_68040 n_72200_68040 Rseg
X1266 n_72200_68040 n_72960_68040 Rseg
X1267 n_72960_68040 n_73340_68040 Rseg
X1268 n_73340_68040 n_73720_68040 Rseg
X1269 n_73720_68040 n_74100_68040 Rseg
X1270 n_74100_68040 n_74860_68040 Rseg
X1271 n_74860_68040 n_75240_68040 Rseg
X1272 n_75240_68040 n_76000_68040 Rseg
X1273 n_76000_68040 n_76380_68040 Rseg
X1274 n_76380_68040 n_76760_68040 Rseg
X1275 n_76760_68040 n_77140_68040 Rseg
X1276 n_77140_68040 n_77520_68040 Rseg
X1277 n_77520_68040 n_77900_68040 Rseg
X1278 n_77900_68040 n_78280_68040 Rseg
X1279 n_78280_68040 n_78660_68040 Rseg
X1280 n_78660_68040 n_79040_68040 Rseg
X1281 n_79040_68040 n_80180_68040 Rseg
X1282 n_80180_68040 n_80560_68040 Rseg
X1283 n_80560_68040 n_80940_68040 Rseg
X1284 n_80940_68040 n_81700_68040 Rseg
X1285 n_81700_68040 n_82080_68040 Rseg
X1286 n_82080_68040 n_83220_68040 Rseg
X1287 n_83220_68040 n_83600_68040 Rseg
X1288 n_83600_68040 n_84740_68040 Rseg
X1289 n_84740_68040 n_85120_68040 Rseg
X1290 n_85120_68040 n_85500_68040 Rseg
X1291 n_85500_68040 n_85880_68040 Rseg
X1292 n_85880_68040 n_86260_68040 Rseg
X1293 n_86260_68040 n_87020_68040 Rseg
X1294 n_87020_68040 n_87400_68040 Rseg
X1295 n_87400_68040 n_87780_68040 Rseg
X1296 n_87780_68040 n_88160_68040 Rseg
X1297 n_88160_68040 n_88540_68040 Rseg
X1298 n_88540_68040 n_88920_68040 Rseg
X1299 n_88920_68040 n_89300_68040 Rseg
X1300 n_89300_68040 n_90060_68040 Rseg
X1301 n_90060_68040 n_90440_68040 Rseg
X1302 n_90440_68040 n_90820_68040 Rseg
X1303 n_90820_68040 n_91200_68040 Rseg
X1304 n_91200_68040 n_91580_68040 Rseg
X1305 n_91580_68040 n_91960_68040 Rseg
X1306 n_91960_68040 n_92340_68040 Rseg
X1307 n_92340_68040 n_92720_68040 Rseg
X1308 n_92720_68040 n_93100_68040 Rseg
X1309 n_93100_68040 n_93480_68040 Rseg
X1310 n_40280_70840 n_40660_70840 Rseg
X1311 n_40660_70840 n_41420_70840 Rseg
X1312 n_41420_70840 n_41800_70840 Rseg
X1313 n_41800_70840 n_42180_70840 Rseg
X1314 n_42180_70840 n_42940_70840 Rseg
X1315 n_42940_70840 n_43320_70840 Rseg
X1316 n_43320_70840 n_43700_70840 Rseg
X1317 n_43700_70840 n_44080_70840 Rseg
X1318 n_44080_70840 n_44460_70840 Rseg
X1319 n_44460_70840 n_44840_70840 Rseg
X1320 n_44840_70840 n_45220_70840 Rseg
X1321 n_45220_70840 n_45600_70840 Rseg
X1322 n_45600_70840 n_46360_70840 Rseg
X1323 n_46360_70840 n_46740_70840 Rseg
X1324 n_46740_70840 n_47120_70840 Rseg
X1325 n_47120_70840 n_47500_70840 Rseg
X1326 n_47500_70840 n_47880_70840 Rseg
X1327 n_47880_70840 n_48260_70840 Rseg
X1328 n_48260_70840 n_48640_70840 Rseg
X1329 n_48640_70840 n_49020_70840 Rseg
X1330 n_49020_70840 n_49400_70840 Rseg
X1331 n_49400_70840 n_49780_70840 Rseg
X1332 n_49780_70840 n_50160_70840 Rseg
X1333 n_50160_70840 n_50540_70840 Rseg
X1334 n_50540_70840 n_50920_70840 Rseg
X1335 n_50920_70840 n_51300_70840 Rseg
X1336 n_51300_70840 n_51680_70840 Rseg
X1337 n_51680_70840 n_52060_70840 Rseg
X1338 n_52060_70840 n_52440_70840 Rseg
X1339 n_52440_70840 n_52820_70840 Rseg
X1340 n_52820_70840 n_53200_70840 Rseg
X1341 n_53200_70840 n_53580_70840 Rseg
X1342 n_53580_70840 n_53960_70840 Rseg
X1343 n_53960_70840 n_54340_70840 Rseg
X1344 n_54340_70840 n_54720_70840 Rseg
X1345 n_54720_70840 n_55100_70840 Rseg
X1346 n_55100_70840 n_55480_70840 Rseg
X1347 n_55480_70840 n_55860_70840 Rseg
X1348 n_55860_70840 n_56240_70840 Rseg
X1349 n_56240_70840 n_56620_70840 Rseg
X1350 n_56620_70840 n_57000_70840 Rseg
X1351 n_57000_70840 n_57380_70840 Rseg
X1352 n_57380_70840 n_57760_70840 Rseg
X1353 n_57760_70840 n_58140_70840 Rseg
X1354 n_58140_70840 n_58520_70840 Rseg
X1355 n_58520_70840 n_58900_70840 Rseg
X1356 n_58900_70840 n_59280_70840 Rseg
X1357 n_59280_70840 n_59660_70840 Rseg
X1358 n_59660_70840 n_60040_70840 Rseg
X1359 n_60040_70840 n_60420_70840 Rseg
X1360 n_60420_70840 n_60800_70840 Rseg
X1361 n_60800_70840 n_61180_70840 Rseg
X1362 n_61180_70840 n_61560_70840 Rseg
X1363 n_61560_70840 n_61940_70840 Rseg
X1364 n_61940_70840 n_62320_70840 Rseg
X1365 n_62320_70840 n_63080_70840 Rseg
X1366 n_63080_70840 n_63460_70840 Rseg
X1367 n_63460_70840 n_63840_70840 Rseg
X1368 n_63840_70840 n_64220_70840 Rseg
X1369 n_64220_70840 n_64600_70840 Rseg
X1370 n_64600_70840 n_64980_70840 Rseg
X1371 n_64980_70840 n_65360_70840 Rseg
X1372 n_65360_70840 n_65740_70840 Rseg
X1373 n_65740_70840 n_66120_70840 Rseg
X1374 n_66120_70840 n_66880_70840 Rseg
X1375 n_66880_70840 n_67260_70840 Rseg
X1376 n_67260_70840 n_68020_70840 Rseg
X1377 n_68020_70840 n_68400_70840 Rseg
X1378 n_68400_70840 n_68780_70840 Rseg
X1379 n_68780_70840 n_69160_70840 Rseg
X1380 n_69160_70840 n_69920_70840 Rseg
X1381 n_69920_70840 n_70300_70840 Rseg
X1382 n_70300_70840 n_71060_70840 Rseg
X1383 n_71060_70840 n_71820_70840 Rseg
X1384 n_71820_70840 n_72200_70840 Rseg
X1385 n_72200_70840 n_72960_70840 Rseg
X1386 n_72960_70840 n_73340_70840 Rseg
X1387 n_73340_70840 n_73720_70840 Rseg
X1388 n_73720_70840 n_74100_70840 Rseg
X1389 n_74100_70840 n_74860_70840 Rseg
X1390 n_74860_70840 n_75240_70840 Rseg
X1391 n_75240_70840 n_76000_70840 Rseg
X1392 n_76000_70840 n_76380_70840 Rseg
X1393 n_76380_70840 n_76760_70840 Rseg
X1394 n_76760_70840 n_77140_70840 Rseg
X1395 n_77140_70840 n_77520_70840 Rseg
X1396 n_77520_70840 n_77900_70840 Rseg
X1397 n_77900_70840 n_78280_70840 Rseg
X1398 n_78280_70840 n_78660_70840 Rseg
X1399 n_78660_70840 n_79040_70840 Rseg
X1400 n_79040_70840 n_80180_70840 Rseg
X1401 n_80180_70840 n_80560_70840 Rseg
X1402 n_80560_70840 n_80940_70840 Rseg
X1403 n_80940_70840 n_81700_70840 Rseg
X1404 n_81700_70840 n_82080_70840 Rseg
X1405 n_82080_70840 n_83220_70840 Rseg
X1406 n_83220_70840 n_83600_70840 Rseg
X1407 n_83600_70840 n_84740_70840 Rseg
X1408 n_84740_70840 n_85120_70840 Rseg
X1409 n_85120_70840 n_85500_70840 Rseg
X1410 n_85500_70840 n_85880_70840 Rseg
X1411 n_85880_70840 n_86260_70840 Rseg
X1412 n_86260_70840 n_87020_70840 Rseg
X1413 n_87020_70840 n_87400_70840 Rseg
X1414 n_87400_70840 n_87780_70840 Rseg
X1415 n_87780_70840 n_88160_70840 Rseg
X1416 n_88160_70840 n_88540_70840 Rseg
X1417 n_88540_70840 n_88920_70840 Rseg
X1418 n_88920_70840 n_89300_70840 Rseg
X1419 n_89300_70840 n_90060_70840 Rseg
X1420 n_90060_70840 n_90440_70840 Rseg
X1421 n_90440_70840 n_90820_70840 Rseg
X1422 n_90820_70840 n_91200_70840 Rseg
X1423 n_91200_70840 n_91580_70840 Rseg
X1424 n_91580_70840 n_91960_70840 Rseg
X1425 n_91960_70840 n_92340_70840 Rseg
X1426 n_92340_70840 n_92720_70840 Rseg
X1427 n_92720_70840 n_93100_70840 Rseg
X1428 n_93100_70840 n_93480_70840 Rseg
X1429 n_40280_73640 n_40660_73640 Rseg
X1430 n_40660_73640 n_41420_73640 Rseg
X1431 n_41420_73640 n_41800_73640 Rseg
X1432 n_41800_73640 n_42180_73640 Rseg
X1433 n_42180_73640 n_42940_73640 Rseg
X1434 n_42940_73640 n_43320_73640 Rseg
X1435 n_43320_73640 n_43700_73640 Rseg
X1436 n_43700_73640 n_44080_73640 Rseg
X1437 n_44080_73640 n_44460_73640 Rseg
X1438 n_44460_73640 n_44840_73640 Rseg
X1439 n_44840_73640 n_45220_73640 Rseg
X1440 n_45220_73640 n_45600_73640 Rseg
X1441 n_45600_73640 n_46360_73640 Rseg
X1442 n_46360_73640 n_46740_73640 Rseg
X1443 n_46740_73640 n_47120_73640 Rseg
X1444 n_47120_73640 n_47500_73640 Rseg
X1445 n_47500_73640 n_47880_73640 Rseg
X1446 n_47880_73640 n_48260_73640 Rseg
X1447 n_48260_73640 n_48640_73640 Rseg
X1448 n_48640_73640 n_49020_73640 Rseg
X1449 n_49020_73640 n_49400_73640 Rseg
X1450 n_49400_73640 n_49780_73640 Rseg
X1451 n_49780_73640 n_50160_73640 Rseg
X1452 n_50160_73640 n_50540_73640 Rseg
X1453 n_50540_73640 n_50920_73640 Rseg
X1454 n_50920_73640 n_51300_73640 Rseg
X1455 n_51300_73640 n_51680_73640 Rseg
X1456 n_51680_73640 n_52060_73640 Rseg
X1457 n_52060_73640 n_52440_73640 Rseg
X1458 n_52440_73640 n_52820_73640 Rseg
X1459 n_52820_73640 n_53200_73640 Rseg
X1460 n_53200_73640 n_53580_73640 Rseg
X1461 n_53580_73640 n_53960_73640 Rseg
X1462 n_53960_73640 n_54340_73640 Rseg
X1463 n_54340_73640 n_54720_73640 Rseg
X1464 n_54720_73640 n_55100_73640 Rseg
X1465 n_55100_73640 n_55480_73640 Rseg
X1466 n_55480_73640 n_55860_73640 Rseg
X1467 n_55860_73640 n_56240_73640 Rseg
X1468 n_56240_73640 n_56620_73640 Rseg
X1469 n_56620_73640 n_57000_73640 Rseg
X1470 n_57000_73640 n_57380_73640 Rseg
X1471 n_57380_73640 n_57760_73640 Rseg
X1472 n_57760_73640 n_58140_73640 Rseg
X1473 n_58140_73640 n_58520_73640 Rseg
X1474 n_58520_73640 n_58900_73640 Rseg
X1475 n_58900_73640 n_59280_73640 Rseg
X1476 n_59280_73640 n_59660_73640 Rseg
X1477 n_59660_73640 n_60040_73640 Rseg
X1478 n_60040_73640 n_60420_73640 Rseg
X1479 n_60420_73640 n_60800_73640 Rseg
X1480 n_60800_73640 n_61180_73640 Rseg
X1481 n_61180_73640 n_61560_73640 Rseg
X1482 n_61560_73640 n_61940_73640 Rseg
X1483 n_61940_73640 n_62320_73640 Rseg
X1484 n_62320_73640 n_63080_73640 Rseg
X1485 n_63080_73640 n_63460_73640 Rseg
X1486 n_63460_73640 n_63840_73640 Rseg
X1487 n_63840_73640 n_64220_73640 Rseg
X1488 n_64220_73640 n_64600_73640 Rseg
X1489 n_64600_73640 n_64980_73640 Rseg
X1490 n_64980_73640 n_65360_73640 Rseg
X1491 n_65360_73640 n_65740_73640 Rseg
X1492 n_65740_73640 n_66120_73640 Rseg
X1493 n_66120_73640 n_66880_73640 Rseg
X1494 n_66880_73640 n_67260_73640 Rseg
X1495 n_67260_73640 n_68020_73640 Rseg
X1496 n_68020_73640 n_68400_73640 Rseg
X1497 n_68400_73640 n_68780_73640 Rseg
X1498 n_68780_73640 n_69160_73640 Rseg
X1499 n_69160_73640 n_69920_73640 Rseg
X1500 n_69920_73640 n_70300_73640 Rseg
X1501 n_70300_73640 n_71060_73640 Rseg
X1502 n_71060_73640 n_71820_73640 Rseg
X1503 n_71820_73640 n_72200_73640 Rseg
X1504 n_72200_73640 n_72960_73640 Rseg
X1505 n_72960_73640 n_73340_73640 Rseg
X1506 n_73340_73640 n_73720_73640 Rseg
X1507 n_73720_73640 n_74100_73640 Rseg
X1508 n_74100_73640 n_74860_73640 Rseg
X1509 n_74860_73640 n_75240_73640 Rseg
X1510 n_75240_73640 n_76000_73640 Rseg
X1511 n_76000_73640 n_76380_73640 Rseg
X1512 n_76380_73640 n_76760_73640 Rseg
X1513 n_76760_73640 n_77140_73640 Rseg
X1514 n_77140_73640 n_77520_73640 Rseg
X1515 n_77520_73640 n_77900_73640 Rseg
X1516 n_77900_73640 n_78280_73640 Rseg
X1517 n_78280_73640 n_78660_73640 Rseg
X1518 n_78660_73640 n_79040_73640 Rseg
X1519 n_79040_73640 n_80180_73640 Rseg
X1520 n_80180_73640 n_80560_73640 Rseg
X1521 n_80560_73640 n_80940_73640 Rseg
X1522 n_80940_73640 n_81700_73640 Rseg
X1523 n_81700_73640 n_82080_73640 Rseg
X1524 n_82080_73640 n_83220_73640 Rseg
X1525 n_83220_73640 n_83600_73640 Rseg
X1526 n_83600_73640 n_84740_73640 Rseg
X1527 n_84740_73640 n_85120_73640 Rseg
X1528 n_85120_73640 n_85500_73640 Rseg
X1529 n_85500_73640 n_85880_73640 Rseg
X1530 n_85880_73640 n_86260_73640 Rseg
X1531 n_86260_73640 n_87020_73640 Rseg
X1532 n_87020_73640 n_87400_73640 Rseg
X1533 n_87400_73640 n_87780_73640 Rseg
X1534 n_87780_73640 n_88160_73640 Rseg
X1535 n_88160_73640 n_88540_73640 Rseg
X1536 n_88540_73640 n_88920_73640 Rseg
X1537 n_88920_73640 n_89300_73640 Rseg
X1538 n_89300_73640 n_90060_73640 Rseg
X1539 n_90060_73640 n_90440_73640 Rseg
X1540 n_90440_73640 n_90820_73640 Rseg
X1541 n_90820_73640 n_91200_73640 Rseg
X1542 n_91200_73640 n_91580_73640 Rseg
X1543 n_91580_73640 n_91960_73640 Rseg
X1544 n_91960_73640 n_92340_73640 Rseg
X1545 n_92340_73640 n_92720_73640 Rseg
X1546 n_92720_73640 n_93100_73640 Rseg
X1547 n_93100_73640 n_93480_73640 Rseg
X1548 n_40280_76440 n_40660_76440 Rseg
X1549 n_40660_76440 n_41420_76440 Rseg
X1550 n_41420_76440 n_41800_76440 Rseg
X1551 n_41800_76440 n_42180_76440 Rseg
X1552 n_42180_76440 n_42940_76440 Rseg
X1553 n_42940_76440 n_43320_76440 Rseg
X1554 n_43320_76440 n_43700_76440 Rseg
X1555 n_43700_76440 n_44080_76440 Rseg
X1556 n_44080_76440 n_44460_76440 Rseg
X1557 n_44460_76440 n_44840_76440 Rseg
X1558 n_44840_76440 n_45220_76440 Rseg
X1559 n_45220_76440 n_45600_76440 Rseg
X1560 n_45600_76440 n_46360_76440 Rseg
X1561 n_46360_76440 n_46740_76440 Rseg
X1562 n_46740_76440 n_47120_76440 Rseg
X1563 n_47120_76440 n_47500_76440 Rseg
X1564 n_47500_76440 n_47880_76440 Rseg
X1565 n_47880_76440 n_48260_76440 Rseg
X1566 n_48260_76440 n_48640_76440 Rseg
X1567 n_48640_76440 n_49020_76440 Rseg
X1568 n_49020_76440 n_49400_76440 Rseg
X1569 n_49400_76440 n_49780_76440 Rseg
X1570 n_49780_76440 n_50160_76440 Rseg
X1571 n_50160_76440 n_50540_76440 Rseg
X1572 n_50540_76440 n_50920_76440 Rseg
X1573 n_50920_76440 n_51300_76440 Rseg
X1574 n_51300_76440 n_51680_76440 Rseg
X1575 n_51680_76440 n_52060_76440 Rseg
X1576 n_52060_76440 n_52440_76440 Rseg
X1577 n_52440_76440 n_52820_76440 Rseg
X1578 n_52820_76440 n_53200_76440 Rseg
X1579 n_53200_76440 n_53580_76440 Rseg
X1580 n_53580_76440 n_53960_76440 Rseg
X1581 n_53960_76440 n_54340_76440 Rseg
X1582 n_54340_76440 n_54720_76440 Rseg
X1583 n_54720_76440 n_55100_76440 Rseg
X1584 n_55100_76440 n_55480_76440 Rseg
X1585 n_55480_76440 n_55860_76440 Rseg
X1586 n_55860_76440 n_56240_76440 Rseg
X1587 n_56240_76440 n_56620_76440 Rseg
X1588 n_56620_76440 n_57000_76440 Rseg
X1589 n_57000_76440 n_57380_76440 Rseg
X1590 n_57380_76440 n_57760_76440 Rseg
X1591 n_57760_76440 n_58140_76440 Rseg
X1592 n_58140_76440 n_58520_76440 Rseg
X1593 n_58520_76440 n_58900_76440 Rseg
X1594 n_58900_76440 n_59280_76440 Rseg
X1595 n_59280_76440 n_59660_76440 Rseg
X1596 n_59660_76440 n_60040_76440 Rseg
X1597 n_60040_76440 n_60420_76440 Rseg
X1598 n_60420_76440 n_60800_76440 Rseg
X1599 n_60800_76440 n_61180_76440 Rseg
X1600 n_61180_76440 n_61560_76440 Rseg
X1601 n_61560_76440 n_61940_76440 Rseg
X1602 n_61940_76440 n_62320_76440 Rseg
X1603 n_62320_76440 n_63080_76440 Rseg
X1604 n_63080_76440 n_63460_76440 Rseg
X1605 n_63460_76440 n_63840_76440 Rseg
X1606 n_63840_76440 n_64220_76440 Rseg
X1607 n_64220_76440 n_64600_76440 Rseg
X1608 n_64600_76440 n_64980_76440 Rseg
X1609 n_64980_76440 n_65360_76440 Rseg
X1610 n_65360_76440 n_65740_76440 Rseg
X1611 n_65740_76440 n_66120_76440 Rseg
X1612 n_66120_76440 n_66880_76440 Rseg
X1613 n_66880_76440 n_67260_76440 Rseg
X1614 n_67260_76440 n_68020_76440 Rseg
X1615 n_68020_76440 n_68400_76440 Rseg
X1616 n_68400_76440 n_68780_76440 Rseg
X1617 n_68780_76440 n_69160_76440 Rseg
X1618 n_69160_76440 n_69920_76440 Rseg
X1619 n_69920_76440 n_70300_76440 Rseg
X1620 n_70300_76440 n_71060_76440 Rseg
X1621 n_71060_76440 n_71820_76440 Rseg
X1622 n_71820_76440 n_72200_76440 Rseg
X1623 n_72200_76440 n_72960_76440 Rseg
X1624 n_72960_76440 n_73340_76440 Rseg
X1625 n_73340_76440 n_73720_76440 Rseg
X1626 n_73720_76440 n_74100_76440 Rseg
X1627 n_74100_76440 n_74860_76440 Rseg
X1628 n_74860_76440 n_75240_76440 Rseg
X1629 n_75240_76440 n_76000_76440 Rseg
X1630 n_76000_76440 n_76380_76440 Rseg
X1631 n_76380_76440 n_76760_76440 Rseg
X1632 n_76760_76440 n_77140_76440 Rseg
X1633 n_77140_76440 n_77520_76440 Rseg
X1634 n_77520_76440 n_77900_76440 Rseg
X1635 n_77900_76440 n_78280_76440 Rseg
X1636 n_78280_76440 n_78660_76440 Rseg
X1637 n_78660_76440 n_79040_76440 Rseg
X1638 n_79040_76440 n_80180_76440 Rseg
X1639 n_80180_76440 n_80560_76440 Rseg
X1640 n_80560_76440 n_80940_76440 Rseg
X1641 n_80940_76440 n_81700_76440 Rseg
X1642 n_81700_76440 n_82080_76440 Rseg
X1643 n_82080_76440 n_83220_76440 Rseg
X1644 n_83220_76440 n_83600_76440 Rseg
X1645 n_83600_76440 n_84740_76440 Rseg
X1646 n_84740_76440 n_85120_76440 Rseg
X1647 n_85120_76440 n_85500_76440 Rseg
X1648 n_85500_76440 n_85880_76440 Rseg
X1649 n_85880_76440 n_86260_76440 Rseg
X1650 n_86260_76440 n_87020_76440 Rseg
X1651 n_87020_76440 n_87400_76440 Rseg
X1652 n_87400_76440 n_87780_76440 Rseg
X1653 n_87780_76440 n_88160_76440 Rseg
X1654 n_88160_76440 n_88540_76440 Rseg
X1655 n_88540_76440 n_88920_76440 Rseg
X1656 n_88920_76440 n_89300_76440 Rseg
X1657 n_89300_76440 n_90060_76440 Rseg
X1658 n_90060_76440 n_90440_76440 Rseg
X1659 n_90440_76440 n_90820_76440 Rseg
X1660 n_90820_76440 n_91200_76440 Rseg
X1661 n_91200_76440 n_91580_76440 Rseg
X1662 n_91580_76440 n_91960_76440 Rseg
X1663 n_91960_76440 n_92340_76440 Rseg
X1664 n_92340_76440 n_92720_76440 Rseg
X1665 n_92720_76440 n_93100_76440 Rseg
X1666 n_93100_76440 n_93480_76440 Rseg
X1667 n_40280_79240 n_40660_79240 Rseg
X1668 n_40660_79240 n_41420_79240 Rseg
X1669 n_41420_79240 n_41800_79240 Rseg
X1670 n_41800_79240 n_42180_79240 Rseg
X1671 n_42180_79240 n_42940_79240 Rseg
X1672 n_42940_79240 n_43320_79240 Rseg
X1673 n_43320_79240 n_43700_79240 Rseg
X1674 n_43700_79240 n_44080_79240 Rseg
X1675 n_44080_79240 n_44460_79240 Rseg
X1676 n_44460_79240 n_44840_79240 Rseg
X1677 n_44840_79240 n_45220_79240 Rseg
X1678 n_45220_79240 n_45600_79240 Rseg
X1679 n_45600_79240 n_46360_79240 Rseg
X1680 n_46360_79240 n_46740_79240 Rseg
X1681 n_46740_79240 n_47120_79240 Rseg
X1682 n_47120_79240 n_47500_79240 Rseg
X1683 n_47500_79240 n_47880_79240 Rseg
X1684 n_47880_79240 n_48260_79240 Rseg
X1685 n_48260_79240 n_48640_79240 Rseg
X1686 n_48640_79240 n_49020_79240 Rseg
X1687 n_49020_79240 n_49400_79240 Rseg
X1688 n_49400_79240 n_49780_79240 Rseg
X1689 n_49780_79240 n_50160_79240 Rseg
X1690 n_50160_79240 n_50540_79240 Rseg
X1691 n_50540_79240 n_50920_79240 Rseg
X1692 n_50920_79240 n_51300_79240 Rseg
X1693 n_51300_79240 n_51680_79240 Rseg
X1694 n_51680_79240 n_52060_79240 Rseg
X1695 n_52060_79240 n_52440_79240 Rseg
X1696 n_52440_79240 n_52820_79240 Rseg
X1697 n_52820_79240 n_53200_79240 Rseg
X1698 n_53200_79240 n_53580_79240 Rseg
X1699 n_53580_79240 n_53960_79240 Rseg
X1700 n_53960_79240 n_54340_79240 Rseg
X1701 n_54340_79240 n_54720_79240 Rseg
X1702 n_54720_79240 n_55100_79240 Rseg
X1703 n_55100_79240 n_55480_79240 Rseg
X1704 n_55480_79240 n_55860_79240 Rseg
X1705 n_55860_79240 n_56240_79240 Rseg
X1706 n_56240_79240 n_56620_79240 Rseg
X1707 n_56620_79240 n_57000_79240 Rseg
X1708 n_57000_79240 n_57380_79240 Rseg
X1709 n_57380_79240 n_57760_79240 Rseg
X1710 n_57760_79240 n_58140_79240 Rseg
X1711 n_58140_79240 n_58520_79240 Rseg
X1712 n_58520_79240 n_58900_79240 Rseg
X1713 n_58900_79240 n_59280_79240 Rseg
X1714 n_59280_79240 n_59660_79240 Rseg
X1715 n_59660_79240 n_60040_79240 Rseg
X1716 n_60040_79240 n_60420_79240 Rseg
X1717 n_60420_79240 n_60800_79240 Rseg
X1718 n_60800_79240 n_61180_79240 Rseg
X1719 n_61180_79240 n_61560_79240 Rseg
X1720 n_61560_79240 n_61940_79240 Rseg
X1721 n_61940_79240 n_62320_79240 Rseg
X1722 n_62320_79240 n_63080_79240 Rseg
X1723 n_63080_79240 n_63460_79240 Rseg
X1724 n_63460_79240 n_63840_79240 Rseg
X1725 n_63840_79240 n_64220_79240 Rseg
X1726 n_64220_79240 n_64600_79240 Rseg
X1727 n_64600_79240 n_64980_79240 Rseg
X1728 n_64980_79240 n_65360_79240 Rseg
X1729 n_65360_79240 n_65740_79240 Rseg
X1730 n_65740_79240 n_66120_79240 Rseg
X1731 n_66120_79240 n_66880_79240 Rseg
X1732 n_66880_79240 n_67260_79240 Rseg
X1733 n_67260_79240 n_68020_79240 Rseg
X1734 n_68020_79240 n_68400_79240 Rseg
X1735 n_68400_79240 n_68780_79240 Rseg
X1736 n_68780_79240 n_69160_79240 Rseg
X1737 n_69160_79240 n_69920_79240 Rseg
X1738 n_69920_79240 n_70300_79240 Rseg
X1739 n_70300_79240 n_71060_79240 Rseg
X1740 n_71060_79240 n_71820_79240 Rseg
X1741 n_71820_79240 n_72200_79240 Rseg
X1742 n_72200_79240 n_72960_79240 Rseg
X1743 n_72960_79240 n_73340_79240 Rseg
X1744 n_73340_79240 n_73720_79240 Rseg
X1745 n_73720_79240 n_74100_79240 Rseg
X1746 n_74100_79240 n_74860_79240 Rseg
X1747 n_74860_79240 n_75240_79240 Rseg
X1748 n_75240_79240 n_76000_79240 Rseg
X1749 n_76000_79240 n_76380_79240 Rseg
X1750 n_76380_79240 n_76760_79240 Rseg
X1751 n_76760_79240 n_77140_79240 Rseg
X1752 n_77140_79240 n_77520_79240 Rseg
X1753 n_77520_79240 n_77900_79240 Rseg
X1754 n_77900_79240 n_78280_79240 Rseg
X1755 n_78280_79240 n_78660_79240 Rseg
X1756 n_78660_79240 n_79040_79240 Rseg
X1757 n_79040_79240 n_80180_79240 Rseg
X1758 n_80180_79240 n_80560_79240 Rseg
X1759 n_80560_79240 n_80940_79240 Rseg
X1760 n_80940_79240 n_81700_79240 Rseg
X1761 n_81700_79240 n_82080_79240 Rseg
X1762 n_82080_79240 n_83220_79240 Rseg
X1763 n_83220_79240 n_83600_79240 Rseg
X1764 n_83600_79240 n_84740_79240 Rseg
X1765 n_84740_79240 n_85120_79240 Rseg
X1766 n_85120_79240 n_85500_79240 Rseg
X1767 n_85500_79240 n_85880_79240 Rseg
X1768 n_85880_79240 n_86260_79240 Rseg
X1769 n_86260_79240 n_87020_79240 Rseg
X1770 n_87020_79240 n_87400_79240 Rseg
X1771 n_87400_79240 n_87780_79240 Rseg
X1772 n_87780_79240 n_88160_79240 Rseg
X1773 n_88160_79240 n_88540_79240 Rseg
X1774 n_88540_79240 n_88920_79240 Rseg
X1775 n_88920_79240 n_89300_79240 Rseg
X1776 n_89300_79240 n_90060_79240 Rseg
X1777 n_90060_79240 n_90440_79240 Rseg
X1778 n_90440_79240 n_90820_79240 Rseg
X1779 n_90820_79240 n_91200_79240 Rseg
X1780 n_91200_79240 n_91580_79240 Rseg
X1781 n_91580_79240 n_91960_79240 Rseg
X1782 n_91960_79240 n_92340_79240 Rseg
X1783 n_92340_79240 n_92720_79240 Rseg
X1784 n_92720_79240 n_93100_79240 Rseg
X1785 n_93100_79240 n_93480_79240 Rseg
X1786 n_40280_82040 n_40660_82040 Rseg
X1787 n_40660_82040 n_41420_82040 Rseg
X1788 n_41420_82040 n_41800_82040 Rseg
X1789 n_41800_82040 n_42180_82040 Rseg
X1790 n_42180_82040 n_42940_82040 Rseg
X1791 n_42940_82040 n_43320_82040 Rseg
X1792 n_43320_82040 n_43700_82040 Rseg
X1793 n_43700_82040 n_44080_82040 Rseg
X1794 n_44080_82040 n_44460_82040 Rseg
X1795 n_44460_82040 n_44840_82040 Rseg
X1796 n_44840_82040 n_45220_82040 Rseg
X1797 n_45220_82040 n_45600_82040 Rseg
X1798 n_45600_82040 n_46360_82040 Rseg
X1799 n_46360_82040 n_46740_82040 Rseg
X1800 n_46740_82040 n_47120_82040 Rseg
X1801 n_47120_82040 n_47500_82040 Rseg
X1802 n_47500_82040 n_47880_82040 Rseg
X1803 n_47880_82040 n_48260_82040 Rseg
X1804 n_48260_82040 n_48640_82040 Rseg
X1805 n_48640_82040 n_49020_82040 Rseg
X1806 n_49020_82040 n_49400_82040 Rseg
X1807 n_49400_82040 n_49780_82040 Rseg
X1808 n_49780_82040 n_50160_82040 Rseg
X1809 n_50160_82040 n_50540_82040 Rseg
X1810 n_50540_82040 n_50920_82040 Rseg
X1811 n_50920_82040 n_51300_82040 Rseg
X1812 n_51300_82040 n_51680_82040 Rseg
X1813 n_51680_82040 n_52060_82040 Rseg
X1814 n_52060_82040 n_52440_82040 Rseg
X1815 n_52440_82040 n_52820_82040 Rseg
X1816 n_52820_82040 n_53200_82040 Rseg
X1817 n_53200_82040 n_53580_82040 Rseg
X1818 n_53580_82040 n_53960_82040 Rseg
X1819 n_53960_82040 n_54340_82040 Rseg
X1820 n_54340_82040 n_54720_82040 Rseg
X1821 n_54720_82040 n_55100_82040 Rseg
X1822 n_55100_82040 n_55480_82040 Rseg
X1823 n_55480_82040 n_55860_82040 Rseg
X1824 n_55860_82040 n_56240_82040 Rseg
X1825 n_56240_82040 n_56620_82040 Rseg
X1826 n_56620_82040 n_57000_82040 Rseg
X1827 n_57000_82040 n_57380_82040 Rseg
X1828 n_57380_82040 n_57760_82040 Rseg
X1829 n_57760_82040 n_58140_82040 Rseg
X1830 n_58140_82040 n_58520_82040 Rseg
X1831 n_58520_82040 n_58900_82040 Rseg
X1832 n_58900_82040 n_59280_82040 Rseg
X1833 n_59280_82040 n_59660_82040 Rseg
X1834 n_59660_82040 n_60040_82040 Rseg
X1835 n_60040_82040 n_60420_82040 Rseg
X1836 n_60420_82040 n_60800_82040 Rseg
X1837 n_60800_82040 n_61180_82040 Rseg
X1838 n_61180_82040 n_61560_82040 Rseg
X1839 n_61560_82040 n_61940_82040 Rseg
X1840 n_61940_82040 n_62320_82040 Rseg
X1841 n_62320_82040 n_63080_82040 Rseg
X1842 n_63080_82040 n_63460_82040 Rseg
X1843 n_63460_82040 n_63840_82040 Rseg
X1844 n_63840_82040 n_64220_82040 Rseg
X1845 n_64220_82040 n_64600_82040 Rseg
X1846 n_64600_82040 n_64980_82040 Rseg
X1847 n_64980_82040 n_65360_82040 Rseg
X1848 n_65360_82040 n_65740_82040 Rseg
X1849 n_65740_82040 n_66120_82040 Rseg
X1850 n_66120_82040 n_66880_82040 Rseg
X1851 n_66880_82040 n_67260_82040 Rseg
X1852 n_67260_82040 n_68020_82040 Rseg
X1853 n_68020_82040 n_68400_82040 Rseg
X1854 n_68400_82040 n_68780_82040 Rseg
X1855 n_68780_82040 n_69160_82040 Rseg
X1856 n_69160_82040 n_69920_82040 Rseg
X1857 n_69920_82040 n_70300_82040 Rseg
X1858 n_70300_82040 n_71060_82040 Rseg
X1859 n_71060_82040 n_71820_82040 Rseg
X1860 n_71820_82040 n_72200_82040 Rseg
X1861 n_72200_82040 n_72960_82040 Rseg
X1862 n_72960_82040 n_73340_82040 Rseg
X1863 n_73340_82040 n_73720_82040 Rseg
X1864 n_73720_82040 n_74100_82040 Rseg
X1865 n_74100_82040 n_74860_82040 Rseg
X1866 n_74860_82040 n_75240_82040 Rseg
X1867 n_75240_82040 n_76000_82040 Rseg
X1868 n_76000_82040 n_76380_82040 Rseg
X1869 n_76380_82040 n_76760_82040 Rseg
X1870 n_76760_82040 n_77140_82040 Rseg
X1871 n_77140_82040 n_77520_82040 Rseg
X1872 n_77520_82040 n_77900_82040 Rseg
X1873 n_77900_82040 n_78280_82040 Rseg
X1874 n_78280_82040 n_78660_82040 Rseg
X1875 n_78660_82040 n_79040_82040 Rseg
X1876 n_79040_82040 n_80180_82040 Rseg
X1877 n_80180_82040 n_80560_82040 Rseg
X1878 n_80560_82040 n_80940_82040 Rseg
X1879 n_80940_82040 n_81700_82040 Rseg
X1880 n_81700_82040 n_82080_82040 Rseg
X1881 n_82080_82040 n_83220_82040 Rseg
X1882 n_83220_82040 n_83600_82040 Rseg
X1883 n_83600_82040 n_84740_82040 Rseg
X1884 n_84740_82040 n_85120_82040 Rseg
X1885 n_85120_82040 n_85500_82040 Rseg
X1886 n_85500_82040 n_85880_82040 Rseg
X1887 n_85880_82040 n_86260_82040 Rseg
X1888 n_86260_82040 n_87020_82040 Rseg
X1889 n_87020_82040 n_87400_82040 Rseg
X1890 n_87400_82040 n_87780_82040 Rseg
X1891 n_87780_82040 n_88160_82040 Rseg
X1892 n_88160_82040 n_88540_82040 Rseg
X1893 n_88540_82040 n_88920_82040 Rseg
X1894 n_88920_82040 n_89300_82040 Rseg
X1895 n_89300_82040 n_90060_82040 Rseg
X1896 n_90060_82040 n_90440_82040 Rseg
X1897 n_90440_82040 n_90820_82040 Rseg
X1898 n_90820_82040 n_91200_82040 Rseg
X1899 n_91200_82040 n_91580_82040 Rseg
X1900 n_91580_82040 n_91960_82040 Rseg
X1901 n_91960_82040 n_92340_82040 Rseg
X1902 n_92340_82040 n_92720_82040 Rseg
X1903 n_92720_82040 n_93100_82040 Rseg
X1904 n_93100_82040 n_93480_82040 Rseg
X1905 n_40280_84840 n_40660_84840 Rseg
X1906 n_40660_84840 n_41420_84840 Rseg
X1907 n_41420_84840 n_41800_84840 Rseg
X1908 n_41800_84840 n_42180_84840 Rseg
X1909 n_42180_84840 n_42940_84840 Rseg
X1910 n_42940_84840 n_43320_84840 Rseg
X1911 n_43320_84840 n_43700_84840 Rseg
X1912 n_43700_84840 n_44080_84840 Rseg
X1913 n_44080_84840 n_44460_84840 Rseg
X1914 n_44460_84840 n_44840_84840 Rseg
X1915 n_44840_84840 n_45220_84840 Rseg
X1916 n_45220_84840 n_45600_84840 Rseg
X1917 n_45600_84840 n_46360_84840 Rseg
X1918 n_46360_84840 n_46740_84840 Rseg
X1919 n_46740_84840 n_47120_84840 Rseg
X1920 n_47120_84840 n_47500_84840 Rseg
X1921 n_47500_84840 n_47880_84840 Rseg
X1922 n_47880_84840 n_48260_84840 Rseg
X1923 n_48260_84840 n_48640_84840 Rseg
X1924 n_48640_84840 n_49020_84840 Rseg
X1925 n_49020_84840 n_49400_84840 Rseg
X1926 n_49400_84840 n_49780_84840 Rseg
X1927 n_49780_84840 n_50160_84840 Rseg
X1928 n_50160_84840 n_50540_84840 Rseg
X1929 n_50540_84840 n_50920_84840 Rseg
X1930 n_50920_84840 n_51300_84840 Rseg
X1931 n_51300_84840 n_51680_84840 Rseg
X1932 n_51680_84840 n_52060_84840 Rseg
X1933 n_52060_84840 n_52440_84840 Rseg
X1934 n_52440_84840 n_52820_84840 Rseg
X1935 n_52820_84840 n_53200_84840 Rseg
X1936 n_53200_84840 n_53580_84840 Rseg
X1937 n_53580_84840 n_53960_84840 Rseg
X1938 n_53960_84840 n_54340_84840 Rseg
X1939 n_54340_84840 n_54720_84840 Rseg
X1940 n_54720_84840 n_55100_84840 Rseg
X1941 n_55100_84840 n_55480_84840 Rseg
X1942 n_55480_84840 n_55860_84840 Rseg
X1943 n_55860_84840 n_56240_84840 Rseg
X1944 n_56240_84840 n_56620_84840 Rseg
X1945 n_56620_84840 n_57000_84840 Rseg
X1946 n_57000_84840 n_57380_84840 Rseg
X1947 n_57380_84840 n_57760_84840 Rseg
X1948 n_57760_84840 n_58140_84840 Rseg
X1949 n_58140_84840 n_58520_84840 Rseg
X1950 n_58520_84840 n_58900_84840 Rseg
X1951 n_58900_84840 n_59280_84840 Rseg
X1952 n_59280_84840 n_59660_84840 Rseg
X1953 n_59660_84840 n_60040_84840 Rseg
X1954 n_60040_84840 n_60420_84840 Rseg
X1955 n_60420_84840 n_60800_84840 Rseg
X1956 n_60800_84840 n_61180_84840 Rseg
X1957 n_61180_84840 n_61560_84840 Rseg
X1958 n_61560_84840 n_61940_84840 Rseg
X1959 n_61940_84840 n_62320_84840 Rseg
X1960 n_62320_84840 n_63080_84840 Rseg
X1961 n_63080_84840 n_63460_84840 Rseg
X1962 n_63460_84840 n_63840_84840 Rseg
X1963 n_63840_84840 n_64220_84840 Rseg
X1964 n_64220_84840 n_64600_84840 Rseg
X1965 n_64600_84840 n_64980_84840 Rseg
X1966 n_64980_84840 n_65360_84840 Rseg
X1967 n_65360_84840 n_65740_84840 Rseg
X1968 n_65740_84840 n_66120_84840 Rseg
X1969 n_66120_84840 n_66880_84840 Rseg
X1970 n_66880_84840 n_67260_84840 Rseg
X1971 n_67260_84840 n_68020_84840 Rseg
X1972 n_68020_84840 n_68400_84840 Rseg
X1973 n_68400_84840 n_68780_84840 Rseg
X1974 n_68780_84840 n_69160_84840 Rseg
X1975 n_69160_84840 n_69920_84840 Rseg
X1976 n_69920_84840 n_70300_84840 Rseg
X1977 n_70300_84840 n_71060_84840 Rseg
X1978 n_71060_84840 n_71820_84840 Rseg
X1979 n_71820_84840 n_72200_84840 Rseg
X1980 n_72200_84840 n_72960_84840 Rseg
X1981 n_72960_84840 n_73340_84840 Rseg
X1982 n_73340_84840 n_73720_84840 Rseg
X1983 n_73720_84840 n_74100_84840 Rseg
X1984 n_74100_84840 n_74860_84840 Rseg
X1985 n_74860_84840 n_75240_84840 Rseg
X1986 n_75240_84840 n_76000_84840 Rseg
X1987 n_76000_84840 n_76380_84840 Rseg
X1988 n_76380_84840 n_76760_84840 Rseg
X1989 n_76760_84840 n_77140_84840 Rseg
X1990 n_77140_84840 n_77520_84840 Rseg
X1991 n_77520_84840 n_77900_84840 Rseg
X1992 n_77900_84840 n_78280_84840 Rseg
X1993 n_78280_84840 n_78660_84840 Rseg
X1994 n_78660_84840 n_79040_84840 Rseg
X1995 n_79040_84840 n_80180_84840 Rseg
X1996 n_80180_84840 n_80560_84840 Rseg
X1997 n_80560_84840 n_80940_84840 Rseg
X1998 n_80940_84840 n_81700_84840 Rseg
X1999 n_81700_84840 n_82080_84840 Rseg
X2000 n_82080_84840 n_83220_84840 Rseg
X2001 n_83220_84840 n_83600_84840 Rseg
X2002 n_83600_84840 n_84740_84840 Rseg
X2003 n_84740_84840 n_85120_84840 Rseg
X2004 n_85120_84840 n_85500_84840 Rseg
X2005 n_85500_84840 n_85880_84840 Rseg
X2006 n_85880_84840 n_86260_84840 Rseg
X2007 n_86260_84840 n_87020_84840 Rseg
X2008 n_87020_84840 n_87400_84840 Rseg
X2009 n_87400_84840 n_87780_84840 Rseg
X2010 n_87780_84840 n_88160_84840 Rseg
X2011 n_88160_84840 n_88540_84840 Rseg
X2012 n_88540_84840 n_88920_84840 Rseg
X2013 n_88920_84840 n_89300_84840 Rseg
X2014 n_89300_84840 n_90060_84840 Rseg
X2015 n_90060_84840 n_90440_84840 Rseg
X2016 n_90440_84840 n_90820_84840 Rseg
X2017 n_90820_84840 n_91200_84840 Rseg
X2018 n_91200_84840 n_91580_84840 Rseg
X2019 n_91580_84840 n_91960_84840 Rseg
X2020 n_91960_84840 n_92340_84840 Rseg
X2021 n_92340_84840 n_92720_84840 Rseg
X2022 n_92720_84840 n_93100_84840 Rseg
X2023 n_93100_84840 n_93480_84840 Rseg
X2024 n_40280_87640 n_40660_87640 Rseg
X2025 n_40660_87640 n_41420_87640 Rseg
X2026 n_41420_87640 n_41800_87640 Rseg
X2027 n_41800_87640 n_42180_87640 Rseg
X2028 n_42180_87640 n_42940_87640 Rseg
X2029 n_42940_87640 n_43320_87640 Rseg
X2030 n_43320_87640 n_43700_87640 Rseg
X2031 n_43700_87640 n_44080_87640 Rseg
X2032 n_44080_87640 n_44460_87640 Rseg
X2033 n_44460_87640 n_44840_87640 Rseg
X2034 n_44840_87640 n_45220_87640 Rseg
X2035 n_45220_87640 n_45600_87640 Rseg
X2036 n_45600_87640 n_46360_87640 Rseg
X2037 n_46360_87640 n_46740_87640 Rseg
X2038 n_46740_87640 n_47120_87640 Rseg
X2039 n_47120_87640 n_47500_87640 Rseg
X2040 n_47500_87640 n_47880_87640 Rseg
X2041 n_47880_87640 n_48260_87640 Rseg
X2042 n_48260_87640 n_48640_87640 Rseg
X2043 n_48640_87640 n_49020_87640 Rseg
X2044 n_49020_87640 n_49400_87640 Rseg
X2045 n_49400_87640 n_49780_87640 Rseg
X2046 n_49780_87640 n_50160_87640 Rseg
X2047 n_50160_87640 n_50540_87640 Rseg
X2048 n_50540_87640 n_50920_87640 Rseg
X2049 n_50920_87640 n_51300_87640 Rseg
X2050 n_51300_87640 n_51680_87640 Rseg
X2051 n_51680_87640 n_52060_87640 Rseg
X2052 n_52060_87640 n_52440_87640 Rseg
X2053 n_52440_87640 n_52820_87640 Rseg
X2054 n_52820_87640 n_53200_87640 Rseg
X2055 n_53200_87640 n_53580_87640 Rseg
X2056 n_53580_87640 n_53960_87640 Rseg
X2057 n_53960_87640 n_54340_87640 Rseg
X2058 n_54340_87640 n_54720_87640 Rseg
X2059 n_54720_87640 n_55100_87640 Rseg
X2060 n_55100_87640 n_55480_87640 Rseg
X2061 n_55480_87640 n_55860_87640 Rseg
X2062 n_55860_87640 n_56240_87640 Rseg
X2063 n_56240_87640 n_56620_87640 Rseg
X2064 n_56620_87640 n_57000_87640 Rseg
X2065 n_57000_87640 n_57380_87640 Rseg
X2066 n_57380_87640 n_57760_87640 Rseg
X2067 n_57760_87640 n_58140_87640 Rseg
X2068 n_58140_87640 n_58520_87640 Rseg
X2069 n_58520_87640 n_58900_87640 Rseg
X2070 n_58900_87640 n_59280_87640 Rseg
X2071 n_59280_87640 n_59660_87640 Rseg
X2072 n_59660_87640 n_60040_87640 Rseg
X2073 n_60040_87640 n_60420_87640 Rseg
X2074 n_60420_87640 n_60800_87640 Rseg
X2075 n_60800_87640 n_61180_87640 Rseg
X2076 n_61180_87640 n_61560_87640 Rseg
X2077 n_61560_87640 n_61940_87640 Rseg
X2078 n_61940_87640 n_62320_87640 Rseg
X2079 n_62320_87640 n_63080_87640 Rseg
X2080 n_63080_87640 n_63460_87640 Rseg
X2081 n_63460_87640 n_63840_87640 Rseg
X2082 n_63840_87640 n_64220_87640 Rseg
X2083 n_64220_87640 n_64600_87640 Rseg
X2084 n_64600_87640 n_64980_87640 Rseg
X2085 n_64980_87640 n_65360_87640 Rseg
X2086 n_65360_87640 n_65740_87640 Rseg
X2087 n_65740_87640 n_66120_87640 Rseg
X2088 n_66120_87640 n_66880_87640 Rseg
X2089 n_66880_87640 n_67260_87640 Rseg
X2090 n_67260_87640 n_68020_87640 Rseg
X2091 n_68020_87640 n_68400_87640 Rseg
X2092 n_68400_87640 n_68780_87640 Rseg
X2093 n_68780_87640 n_69160_87640 Rseg
X2094 n_69160_87640 n_69920_87640 Rseg
X2095 n_69920_87640 n_70300_87640 Rseg
X2096 n_70300_87640 n_71060_87640 Rseg
X2097 n_71060_87640 n_71820_87640 Rseg
X2098 n_71820_87640 n_72200_87640 Rseg
X2099 n_72200_87640 n_72960_87640 Rseg
X2100 n_72960_87640 n_73340_87640 Rseg
X2101 n_73340_87640 n_73720_87640 Rseg
X2102 n_73720_87640 n_74100_87640 Rseg
X2103 n_74100_87640 n_74860_87640 Rseg
X2104 n_74860_87640 n_75240_87640 Rseg
X2105 n_75240_87640 n_76000_87640 Rseg
X2106 n_76000_87640 n_76380_87640 Rseg
X2107 n_76380_87640 n_76760_87640 Rseg
X2108 n_76760_87640 n_77140_87640 Rseg
X2109 n_77140_87640 n_77520_87640 Rseg
X2110 n_77520_87640 n_77900_87640 Rseg
X2111 n_77900_87640 n_78280_87640 Rseg
X2112 n_78280_87640 n_78660_87640 Rseg
X2113 n_78660_87640 n_79040_87640 Rseg
X2114 n_79040_87640 n_80180_87640 Rseg
X2115 n_80180_87640 n_80560_87640 Rseg
X2116 n_80560_87640 n_80940_87640 Rseg
X2117 n_80940_87640 n_81700_87640 Rseg
X2118 n_81700_87640 n_82080_87640 Rseg
X2119 n_82080_87640 n_83220_87640 Rseg
X2120 n_83220_87640 n_83600_87640 Rseg
X2121 n_83600_87640 n_84740_87640 Rseg
X2122 n_84740_87640 n_85120_87640 Rseg
X2123 n_85120_87640 n_85500_87640 Rseg
X2124 n_85500_87640 n_85880_87640 Rseg
X2125 n_85880_87640 n_86260_87640 Rseg
X2126 n_86260_87640 n_87020_87640 Rseg
X2127 n_87020_87640 n_87400_87640 Rseg
X2128 n_87400_87640 n_87780_87640 Rseg
X2129 n_87780_87640 n_88160_87640 Rseg
X2130 n_88160_87640 n_88540_87640 Rseg
X2131 n_88540_87640 n_88920_87640 Rseg
X2132 n_88920_87640 n_89300_87640 Rseg
X2133 n_89300_87640 n_90060_87640 Rseg
X2134 n_90060_87640 n_90440_87640 Rseg
X2135 n_90440_87640 n_90820_87640 Rseg
X2136 n_90820_87640 n_91200_87640 Rseg
X2137 n_91200_87640 n_91580_87640 Rseg
X2138 n_91580_87640 n_91960_87640 Rseg
X2139 n_91960_87640 n_92340_87640 Rseg
X2140 n_92340_87640 n_92720_87640 Rseg
X2141 n_92720_87640 n_93100_87640 Rseg
X2142 n_93100_87640 n_93480_87640 Rseg
* the vertical resistors:
X2143 n_40280_40040 n_40280_42840 Rseg
X2144 n_40280_42840 n_40280_45640 Rseg
X2145 n_40280_45640 n_40280_48440 Rseg
X2146 n_40280_48440 n_40280_51240 Rseg
X2147 n_40280_51240 n_40280_54040 Rseg
X2148 n_40280_54040 n_40280_56840 Rseg
X2149 n_40280_56840 n_40280_59640 Rseg
X2150 n_40280_59640 n_40280_62440 Rseg
X2151 n_40280_62440 n_40280_65240 Rseg
X2152 n_40280_65240 n_40280_68040 Rseg
X2153 n_40280_68040 n_40280_70840 Rseg
X2154 n_40280_70840 n_40280_73640 Rseg
X2155 n_40280_73640 n_40280_76440 Rseg
X2156 n_40280_76440 n_40280_79240 Rseg
X2157 n_40280_79240 n_40280_82040 Rseg
X2158 n_40280_82040 n_40280_84840 Rseg
X2159 n_40280_84840 n_40280_87640 Rseg
X2160 n_40660_40040 n_40660_42840 Rseg
X2161 n_40660_42840 n_40660_45640 Rseg
X2162 n_40660_45640 n_40660_48440 Rseg
X2163 n_40660_48440 n_40660_51240 Rseg
X2164 n_40660_51240 n_40660_54040 Rseg
X2165 n_40660_54040 n_40660_56840 Rseg
X2166 n_40660_56840 n_40660_59640 Rseg
X2167 n_40660_59640 n_40660_62440 Rseg
X2168 n_40660_62440 n_40660_65240 Rseg
X2169 n_40660_65240 n_40660_68040 Rseg
X2170 n_40660_68040 n_40660_70840 Rseg
X2171 n_40660_70840 n_40660_73640 Rseg
X2172 n_40660_73640 n_40660_76440 Rseg
X2173 n_40660_76440 n_40660_79240 Rseg
X2174 n_40660_79240 n_40660_82040 Rseg
X2175 n_40660_82040 n_40660_84840 Rseg
X2176 n_40660_84840 n_40660_87640 Rseg
X2177 n_41420_40040 n_41420_42840 Rseg
X2178 n_41420_42840 n_41420_45640 Rseg
X2179 n_41420_45640 n_41420_48440 Rseg
X2180 n_41420_48440 n_41420_51240 Rseg
X2181 n_41420_51240 n_41420_54040 Rseg
X2182 n_41420_54040 n_41420_56840 Rseg
X2183 n_41420_56840 n_41420_59640 Rseg
X2184 n_41420_59640 n_41420_62440 Rseg
X2185 n_41420_62440 n_41420_65240 Rseg
X2186 n_41420_65240 n_41420_68040 Rseg
X2187 n_41420_68040 n_41420_70840 Rseg
X2188 n_41420_70840 n_41420_73640 Rseg
X2189 n_41420_73640 n_41420_76440 Rseg
X2190 n_41420_76440 n_41420_79240 Rseg
X2191 n_41420_79240 n_41420_82040 Rseg
X2192 n_41420_82040 n_41420_84840 Rseg
X2193 n_41420_84840 n_41420_87640 Rseg
X2194 n_41800_40040 n_41800_42840 Rseg
X2195 n_41800_42840 n_41800_45640 Rseg
X2196 n_41800_45640 n_41800_48440 Rseg
X2197 n_41800_48440 n_41800_51240 Rseg
X2198 n_41800_51240 n_41800_54040 Rseg
X2199 n_41800_54040 n_41800_56840 Rseg
X2200 n_41800_56840 n_41800_59640 Rseg
X2201 n_41800_59640 n_41800_62440 Rseg
X2202 n_41800_62440 n_41800_65240 Rseg
X2203 n_41800_65240 n_41800_68040 Rseg
X2204 n_41800_68040 n_41800_70840 Rseg
X2205 n_41800_70840 n_41800_73640 Rseg
X2206 n_41800_73640 n_41800_76440 Rseg
X2207 n_41800_76440 n_41800_79240 Rseg
X2208 n_41800_79240 n_41800_82040 Rseg
X2209 n_41800_82040 n_41800_84840 Rseg
X2210 n_41800_84840 n_41800_87640 Rseg
X2211 n_42180_40040 n_42180_42840 Rseg
X2212 n_42180_42840 n_42180_45640 Rseg
X2213 n_42180_45640 n_42180_48440 Rseg
X2214 n_42180_48440 n_42180_51240 Rseg
X2215 n_42180_51240 n_42180_54040 Rseg
X2216 n_42180_54040 n_42180_56840 Rseg
X2217 n_42180_56840 n_42180_59640 Rseg
X2218 n_42180_59640 n_42180_62440 Rseg
X2219 n_42180_62440 n_42180_65240 Rseg
X2220 n_42180_65240 n_42180_68040 Rseg
X2221 n_42180_68040 n_42180_70840 Rseg
X2222 n_42180_70840 n_42180_73640 Rseg
X2223 n_42180_73640 n_42180_76440 Rseg
X2224 n_42180_76440 n_42180_79240 Rseg
X2225 n_42180_79240 n_42180_82040 Rseg
X2226 n_42180_82040 n_42180_84840 Rseg
X2227 n_42180_84840 n_42180_87640 Rseg
X2228 n_42940_40040 n_42940_42840 Rseg
X2229 n_42940_42840 n_42940_45640 Rseg
X2230 n_42940_45640 n_42940_48440 Rseg
X2231 n_42940_48440 n_42940_51240 Rseg
X2232 n_42940_51240 n_42940_54040 Rseg
X2233 n_42940_54040 n_42940_56840 Rseg
X2234 n_42940_56840 n_42940_59640 Rseg
X2235 n_42940_59640 n_42940_62440 Rseg
X2236 n_42940_62440 n_42940_65240 Rseg
X2237 n_42940_65240 n_42940_68040 Rseg
X2238 n_42940_68040 n_42940_70840 Rseg
X2239 n_42940_70840 n_42940_73640 Rseg
X2240 n_42940_73640 n_42940_76440 Rseg
X2241 n_42940_76440 n_42940_79240 Rseg
X2242 n_42940_79240 n_42940_82040 Rseg
X2243 n_42940_82040 n_42940_84840 Rseg
X2244 n_42940_84840 n_42940_87640 Rseg
X2245 n_43320_40040 n_43320_42840 Rseg
X2246 n_43320_42840 n_43320_45640 Rseg
X2247 n_43320_45640 n_43320_48440 Rseg
X2248 n_43320_48440 n_43320_51240 Rseg
X2249 n_43320_51240 n_43320_54040 Rseg
X2250 n_43320_54040 n_43320_56840 Rseg
X2251 n_43320_56840 n_43320_59640 Rseg
X2252 n_43320_59640 n_43320_62440 Rseg
X2253 n_43320_62440 n_43320_65240 Rseg
X2254 n_43320_65240 n_43320_68040 Rseg
X2255 n_43320_68040 n_43320_70840 Rseg
X2256 n_43320_70840 n_43320_73640 Rseg
X2257 n_43320_73640 n_43320_76440 Rseg
X2258 n_43320_76440 n_43320_79240 Rseg
X2259 n_43320_79240 n_43320_82040 Rseg
X2260 n_43320_82040 n_43320_84840 Rseg
X2261 n_43320_84840 n_43320_87640 Rseg
X2262 n_43700_40040 n_43700_42840 Rseg
X2263 n_43700_42840 n_43700_45640 Rseg
X2264 n_43700_45640 n_43700_48440 Rseg
X2265 n_43700_48440 n_43700_51240 Rseg
X2266 n_43700_51240 n_43700_54040 Rseg
X2267 n_43700_54040 n_43700_56840 Rseg
X2268 n_43700_56840 n_43700_59640 Rseg
X2269 n_43700_59640 n_43700_62440 Rseg
X2270 n_43700_62440 n_43700_65240 Rseg
X2271 n_43700_65240 n_43700_68040 Rseg
X2272 n_43700_68040 n_43700_70840 Rseg
X2273 n_43700_70840 n_43700_73640 Rseg
X2274 n_43700_73640 n_43700_76440 Rseg
X2275 n_43700_76440 n_43700_79240 Rseg
X2276 n_43700_79240 n_43700_82040 Rseg
X2277 n_43700_82040 n_43700_84840 Rseg
X2278 n_43700_84840 n_43700_87640 Rseg
X2279 n_44080_40040 n_44080_42840 Rseg
X2280 n_44080_42840 n_44080_45640 Rseg
X2281 n_44080_45640 n_44080_48440 Rseg
X2282 n_44080_48440 n_44080_51240 Rseg
X2283 n_44080_51240 n_44080_54040 Rseg
X2284 n_44080_54040 n_44080_56840 Rseg
X2285 n_44080_56840 n_44080_59640 Rseg
X2286 n_44080_59640 n_44080_62440 Rseg
X2287 n_44080_62440 n_44080_65240 Rseg
X2288 n_44080_65240 n_44080_68040 Rseg
X2289 n_44080_68040 n_44080_70840 Rseg
X2290 n_44080_70840 n_44080_73640 Rseg
X2291 n_44080_73640 n_44080_76440 Rseg
X2292 n_44080_76440 n_44080_79240 Rseg
X2293 n_44080_79240 n_44080_82040 Rseg
X2294 n_44080_82040 n_44080_84840 Rseg
X2295 n_44080_84840 n_44080_87640 Rseg
X2296 n_44460_40040 n_44460_42840 Rseg
X2297 n_44460_42840 n_44460_45640 Rseg
X2298 n_44460_45640 n_44460_48440 Rseg
X2299 n_44460_48440 n_44460_51240 Rseg
X2300 n_44460_51240 n_44460_54040 Rseg
X2301 n_44460_54040 n_44460_56840 Rseg
X2302 n_44460_56840 n_44460_59640 Rseg
X2303 n_44460_59640 n_44460_62440 Rseg
X2304 n_44460_62440 n_44460_65240 Rseg
X2305 n_44460_65240 n_44460_68040 Rseg
X2306 n_44460_68040 n_44460_70840 Rseg
X2307 n_44460_70840 n_44460_73640 Rseg
X2308 n_44460_73640 n_44460_76440 Rseg
X2309 n_44460_76440 n_44460_79240 Rseg
X2310 n_44460_79240 n_44460_82040 Rseg
X2311 n_44460_82040 n_44460_84840 Rseg
X2312 n_44460_84840 n_44460_87640 Rseg
X2313 n_44840_40040 n_44840_42840 Rseg
X2314 n_44840_42840 n_44840_45640 Rseg
X2315 n_44840_45640 n_44840_48440 Rseg
X2316 n_44840_48440 n_44840_51240 Rseg
X2317 n_44840_51240 n_44840_54040 Rseg
X2318 n_44840_54040 n_44840_56840 Rseg
X2319 n_44840_56840 n_44840_59640 Rseg
X2320 n_44840_59640 n_44840_62440 Rseg
X2321 n_44840_62440 n_44840_65240 Rseg
X2322 n_44840_65240 n_44840_68040 Rseg
X2323 n_44840_68040 n_44840_70840 Rseg
X2324 n_44840_70840 n_44840_73640 Rseg
X2325 n_44840_73640 n_44840_76440 Rseg
X2326 n_44840_76440 n_44840_79240 Rseg
X2327 n_44840_79240 n_44840_82040 Rseg
X2328 n_44840_82040 n_44840_84840 Rseg
X2329 n_44840_84840 n_44840_87640 Rseg
X2330 n_45220_40040 n_45220_42840 Rseg
X2331 n_45220_42840 n_45220_45640 Rseg
X2332 n_45220_45640 n_45220_48440 Rseg
X2333 n_45220_48440 n_45220_51240 Rseg
X2334 n_45220_51240 n_45220_54040 Rseg
X2335 n_45220_54040 n_45220_56840 Rseg
X2336 n_45220_56840 n_45220_59640 Rseg
X2337 n_45220_59640 n_45220_62440 Rseg
X2338 n_45220_62440 n_45220_65240 Rseg
X2339 n_45220_65240 n_45220_68040 Rseg
X2340 n_45220_68040 n_45220_70840 Rseg
X2341 n_45220_70840 n_45220_73640 Rseg
X2342 n_45220_73640 n_45220_76440 Rseg
X2343 n_45220_76440 n_45220_79240 Rseg
X2344 n_45220_79240 n_45220_82040 Rseg
X2345 n_45220_82040 n_45220_84840 Rseg
X2346 n_45220_84840 n_45220_87640 Rseg
X2347 n_45600_40040 n_45600_42840 Rseg
X2348 n_45600_42840 n_45600_45640 Rseg
X2349 n_45600_45640 n_45600_48440 Rseg
X2350 n_45600_48440 n_45600_51240 Rseg
X2351 n_45600_51240 n_45600_54040 Rseg
X2352 n_45600_54040 n_45600_56840 Rseg
X2353 n_45600_56840 n_45600_59640 Rseg
X2354 n_45600_59640 n_45600_62440 Rseg
X2355 n_45600_62440 n_45600_65240 Rseg
X2356 n_45600_65240 n_45600_68040 Rseg
X2357 n_45600_68040 n_45600_70840 Rseg
X2358 n_45600_70840 n_45600_73640 Rseg
X2359 n_45600_73640 n_45600_76440 Rseg
X2360 n_45600_76440 n_45600_79240 Rseg
X2361 n_45600_79240 n_45600_82040 Rseg
X2362 n_45600_82040 n_45600_84840 Rseg
X2363 n_45600_84840 n_45600_87640 Rseg
X2364 n_46360_40040 n_46360_42840 Rseg
X2365 n_46360_42840 n_46360_45640 Rseg
X2366 n_46360_45640 n_46360_48440 Rseg
X2367 n_46360_48440 n_46360_51240 Rseg
X2368 n_46360_51240 n_46360_54040 Rseg
X2369 n_46360_54040 n_46360_56840 Rseg
X2370 n_46360_56840 n_46360_59640 Rseg
X2371 n_46360_59640 n_46360_62440 Rseg
X2372 n_46360_62440 n_46360_65240 Rseg
X2373 n_46360_65240 n_46360_68040 Rseg
X2374 n_46360_68040 n_46360_70840 Rseg
X2375 n_46360_70840 n_46360_73640 Rseg
X2376 n_46360_73640 n_46360_76440 Rseg
X2377 n_46360_76440 n_46360_79240 Rseg
X2378 n_46360_79240 n_46360_82040 Rseg
X2379 n_46360_82040 n_46360_84840 Rseg
X2380 n_46360_84840 n_46360_87640 Rseg
X2381 n_46740_40040 n_46740_42840 Rseg
X2382 n_46740_42840 n_46740_45640 Rseg
X2383 n_46740_45640 n_46740_48440 Rseg
X2384 n_46740_48440 n_46740_51240 Rseg
X2385 n_46740_51240 n_46740_54040 Rseg
X2386 n_46740_54040 n_46740_56840 Rseg
X2387 n_46740_56840 n_46740_59640 Rseg
X2388 n_46740_59640 n_46740_62440 Rseg
X2389 n_46740_62440 n_46740_65240 Rseg
X2390 n_46740_65240 n_46740_68040 Rseg
X2391 n_46740_68040 n_46740_70840 Rseg
X2392 n_46740_70840 n_46740_73640 Rseg
X2393 n_46740_73640 n_46740_76440 Rseg
X2394 n_46740_76440 n_46740_79240 Rseg
X2395 n_46740_79240 n_46740_82040 Rseg
X2396 n_46740_82040 n_46740_84840 Rseg
X2397 n_46740_84840 n_46740_87640 Rseg
X2398 n_47120_40040 n_47120_42840 Rseg
X2399 n_47120_42840 n_47120_45640 Rseg
X2400 n_47120_45640 n_47120_48440 Rseg
X2401 n_47120_48440 n_47120_51240 Rseg
X2402 n_47120_51240 n_47120_54040 Rseg
X2403 n_47120_54040 n_47120_56840 Rseg
X2404 n_47120_56840 n_47120_59640 Rseg
X2405 n_47120_59640 n_47120_62440 Rseg
X2406 n_47120_62440 n_47120_65240 Rseg
X2407 n_47120_65240 n_47120_68040 Rseg
X2408 n_47120_68040 n_47120_70840 Rseg
X2409 n_47120_70840 n_47120_73640 Rseg
X2410 n_47120_73640 n_47120_76440 Rseg
X2411 n_47120_76440 n_47120_79240 Rseg
X2412 n_47120_79240 n_47120_82040 Rseg
X2413 n_47120_82040 n_47120_84840 Rseg
X2414 n_47120_84840 n_47120_87640 Rseg
X2415 n_47500_40040 n_47500_42840 Rseg
X2416 n_47500_42840 n_47500_45640 Rseg
X2417 n_47500_45640 n_47500_48440 Rseg
X2418 n_47500_48440 n_47500_51240 Rseg
X2419 n_47500_51240 n_47500_54040 Rseg
X2420 n_47500_54040 n_47500_56840 Rseg
X2421 n_47500_56840 n_47500_59640 Rseg
X2422 n_47500_59640 n_47500_62440 Rseg
X2423 n_47500_62440 n_47500_65240 Rseg
X2424 n_47500_65240 n_47500_68040 Rseg
X2425 n_47500_68040 n_47500_70840 Rseg
X2426 n_47500_70840 n_47500_73640 Rseg
X2427 n_47500_73640 n_47500_76440 Rseg
X2428 n_47500_76440 n_47500_79240 Rseg
X2429 n_47500_79240 n_47500_82040 Rseg
X2430 n_47500_82040 n_47500_84840 Rseg
X2431 n_47500_84840 n_47500_87640 Rseg
X2432 n_47880_40040 n_47880_42840 Rseg
X2433 n_47880_42840 n_47880_45640 Rseg
X2434 n_47880_45640 n_47880_48440 Rseg
X2435 n_47880_48440 n_47880_51240 Rseg
X2436 n_47880_51240 n_47880_54040 Rseg
X2437 n_47880_54040 n_47880_56840 Rseg
X2438 n_47880_56840 n_47880_59640 Rseg
X2439 n_47880_59640 n_47880_62440 Rseg
X2440 n_47880_62440 n_47880_65240 Rseg
X2441 n_47880_65240 n_47880_68040 Rseg
X2442 n_47880_68040 n_47880_70840 Rseg
X2443 n_47880_70840 n_47880_73640 Rseg
X2444 n_47880_73640 n_47880_76440 Rseg
X2445 n_47880_76440 n_47880_79240 Rseg
X2446 n_47880_79240 n_47880_82040 Rseg
X2447 n_47880_82040 n_47880_84840 Rseg
X2448 n_47880_84840 n_47880_87640 Rseg
X2449 n_48260_40040 n_48260_42840 Rseg
X2450 n_48260_42840 n_48260_45640 Rseg
X2451 n_48260_45640 n_48260_48440 Rseg
X2452 n_48260_48440 n_48260_51240 Rseg
X2453 n_48260_51240 n_48260_54040 Rseg
X2454 n_48260_54040 n_48260_56840 Rseg
X2455 n_48260_56840 n_48260_59640 Rseg
X2456 n_48260_59640 n_48260_62440 Rseg
X2457 n_48260_62440 n_48260_65240 Rseg
X2458 n_48260_65240 n_48260_68040 Rseg
X2459 n_48260_68040 n_48260_70840 Rseg
X2460 n_48260_70840 n_48260_73640 Rseg
X2461 n_48260_73640 n_48260_76440 Rseg
X2462 n_48260_76440 n_48260_79240 Rseg
X2463 n_48260_79240 n_48260_82040 Rseg
X2464 n_48260_82040 n_48260_84840 Rseg
X2465 n_48260_84840 n_48260_87640 Rseg
X2466 n_48640_40040 n_48640_42840 Rseg
X2467 n_48640_42840 n_48640_45640 Rseg
X2468 n_48640_45640 n_48640_48440 Rseg
X2469 n_48640_48440 n_48640_51240 Rseg
X2470 n_48640_51240 n_48640_54040 Rseg
X2471 n_48640_54040 n_48640_56840 Rseg
X2472 n_48640_56840 n_48640_59640 Rseg
X2473 n_48640_59640 n_48640_62440 Rseg
X2474 n_48640_62440 n_48640_65240 Rseg
X2475 n_48640_65240 n_48640_68040 Rseg
X2476 n_48640_68040 n_48640_70840 Rseg
X2477 n_48640_70840 n_48640_73640 Rseg
X2478 n_48640_73640 n_48640_76440 Rseg
X2479 n_48640_76440 n_48640_79240 Rseg
X2480 n_48640_79240 n_48640_82040 Rseg
X2481 n_48640_82040 n_48640_84840 Rseg
X2482 n_48640_84840 n_48640_87640 Rseg
X2483 n_49020_40040 n_49020_42840 Rseg
X2484 n_49020_42840 n_49020_45640 Rseg
X2485 n_49020_45640 n_49020_48440 Rseg
X2486 n_49020_48440 n_49020_51240 Rseg
X2487 n_49020_51240 n_49020_54040 Rseg
X2488 n_49020_54040 n_49020_56840 Rseg
X2489 n_49020_56840 n_49020_59640 Rseg
X2490 n_49020_59640 n_49020_62440 Rseg
X2491 n_49020_62440 n_49020_65240 Rseg
X2492 n_49020_65240 n_49020_68040 Rseg
X2493 n_49020_68040 n_49020_70840 Rseg
X2494 n_49020_70840 n_49020_73640 Rseg
X2495 n_49020_73640 n_49020_76440 Rseg
X2496 n_49020_76440 n_49020_79240 Rseg
X2497 n_49020_79240 n_49020_82040 Rseg
X2498 n_49020_82040 n_49020_84840 Rseg
X2499 n_49020_84840 n_49020_87640 Rseg
X2500 n_49400_40040 n_49400_42840 Rseg
X2501 n_49400_42840 n_49400_45640 Rseg
X2502 n_49400_45640 n_49400_48440 Rseg
X2503 n_49400_48440 n_49400_51240 Rseg
X2504 n_49400_51240 n_49400_54040 Rseg
X2505 n_49400_54040 n_49400_56840 Rseg
X2506 n_49400_56840 n_49400_59640 Rseg
X2507 n_49400_59640 n_49400_62440 Rseg
X2508 n_49400_62440 n_49400_65240 Rseg
X2509 n_49400_65240 n_49400_68040 Rseg
X2510 n_49400_68040 n_49400_70840 Rseg
X2511 n_49400_70840 n_49400_73640 Rseg
X2512 n_49400_73640 n_49400_76440 Rseg
X2513 n_49400_76440 n_49400_79240 Rseg
X2514 n_49400_79240 n_49400_82040 Rseg
X2515 n_49400_82040 n_49400_84840 Rseg
X2516 n_49400_84840 n_49400_87640 Rseg
X2517 n_49780_40040 n_49780_42840 Rseg
X2518 n_49780_42840 n_49780_45640 Rseg
X2519 n_49780_45640 n_49780_48440 Rseg
X2520 n_49780_48440 n_49780_51240 Rseg
X2521 n_49780_51240 n_49780_54040 Rseg
X2522 n_49780_54040 n_49780_56840 Rseg
X2523 n_49780_56840 n_49780_59640 Rseg
X2524 n_49780_59640 n_49780_62440 Rseg
X2525 n_49780_62440 n_49780_65240 Rseg
X2526 n_49780_65240 n_49780_68040 Rseg
X2527 n_49780_68040 n_49780_70840 Rseg
X2528 n_49780_70840 n_49780_73640 Rseg
X2529 n_49780_73640 n_49780_76440 Rseg
X2530 n_49780_76440 n_49780_79240 Rseg
X2531 n_49780_79240 n_49780_82040 Rseg
X2532 n_49780_82040 n_49780_84840 Rseg
X2533 n_49780_84840 n_49780_87640 Rseg
X2534 n_50160_40040 n_50160_42840 Rseg
X2535 n_50160_42840 n_50160_45640 Rseg
X2536 n_50160_45640 n_50160_48440 Rseg
X2537 n_50160_48440 n_50160_51240 Rseg
X2538 n_50160_51240 n_50160_54040 Rseg
X2539 n_50160_54040 n_50160_56840 Rseg
X2540 n_50160_56840 n_50160_59640 Rseg
X2541 n_50160_59640 n_50160_62440 Rseg
X2542 n_50160_62440 n_50160_65240 Rseg
X2543 n_50160_65240 n_50160_68040 Rseg
X2544 n_50160_68040 n_50160_70840 Rseg
X2545 n_50160_70840 n_50160_73640 Rseg
X2546 n_50160_73640 n_50160_76440 Rseg
X2547 n_50160_76440 n_50160_79240 Rseg
X2548 n_50160_79240 n_50160_82040 Rseg
X2549 n_50160_82040 n_50160_84840 Rseg
X2550 n_50160_84840 n_50160_87640 Rseg
X2551 n_50540_40040 n_50540_42840 Rseg
X2552 n_50540_42840 n_50540_45640 Rseg
X2553 n_50540_45640 n_50540_48440 Rseg
X2554 n_50540_48440 n_50540_51240 Rseg
X2555 n_50540_51240 n_50540_54040 Rseg
X2556 n_50540_54040 n_50540_56840 Rseg
X2557 n_50540_56840 n_50540_59640 Rseg
X2558 n_50540_59640 n_50540_62440 Rseg
X2559 n_50540_62440 n_50540_65240 Rseg
X2560 n_50540_65240 n_50540_68040 Rseg
X2561 n_50540_68040 n_50540_70840 Rseg
X2562 n_50540_70840 n_50540_73640 Rseg
X2563 n_50540_73640 n_50540_76440 Rseg
X2564 n_50540_76440 n_50540_79240 Rseg
X2565 n_50540_79240 n_50540_82040 Rseg
X2566 n_50540_82040 n_50540_84840 Rseg
X2567 n_50540_84840 n_50540_87640 Rseg
X2568 n_50920_40040 n_50920_42840 Rseg
X2569 n_50920_42840 n_50920_45640 Rseg
X2570 n_50920_45640 n_50920_48440 Rseg
X2571 n_50920_48440 n_50920_51240 Rseg
X2572 n_50920_51240 n_50920_54040 Rseg
X2573 n_50920_54040 n_50920_56840 Rseg
X2574 n_50920_56840 n_50920_59640 Rseg
X2575 n_50920_59640 n_50920_62440 Rseg
X2576 n_50920_62440 n_50920_65240 Rseg
X2577 n_50920_65240 n_50920_68040 Rseg
X2578 n_50920_68040 n_50920_70840 Rseg
X2579 n_50920_70840 n_50920_73640 Rseg
X2580 n_50920_73640 n_50920_76440 Rseg
X2581 n_50920_76440 n_50920_79240 Rseg
X2582 n_50920_79240 n_50920_82040 Rseg
X2583 n_50920_82040 n_50920_84840 Rseg
X2584 n_50920_84840 n_50920_87640 Rseg
X2585 n_51300_40040 n_51300_42840 Rseg
X2586 n_51300_42840 n_51300_45640 Rseg
X2587 n_51300_45640 n_51300_48440 Rseg
X2588 n_51300_48440 n_51300_51240 Rseg
X2589 n_51300_51240 n_51300_54040 Rseg
X2590 n_51300_54040 n_51300_56840 Rseg
X2591 n_51300_56840 n_51300_59640 Rseg
X2592 n_51300_59640 n_51300_62440 Rseg
X2593 n_51300_62440 n_51300_65240 Rseg
X2594 n_51300_65240 n_51300_68040 Rseg
X2595 n_51300_68040 n_51300_70840 Rseg
X2596 n_51300_70840 n_51300_73640 Rseg
X2597 n_51300_73640 n_51300_76440 Rseg
X2598 n_51300_76440 n_51300_79240 Rseg
X2599 n_51300_79240 n_51300_82040 Rseg
X2600 n_51300_82040 n_51300_84840 Rseg
X2601 n_51300_84840 n_51300_87640 Rseg
X2602 n_51680_40040 n_51680_42840 Rseg
X2603 n_51680_42840 n_51680_45640 Rseg
X2604 n_51680_45640 n_51680_48440 Rseg
X2605 n_51680_48440 n_51680_51240 Rseg
X2606 n_51680_51240 n_51680_54040 Rseg
X2607 n_51680_54040 n_51680_56840 Rseg
X2608 n_51680_56840 n_51680_59640 Rseg
X2609 n_51680_59640 n_51680_62440 Rseg
X2610 n_51680_62440 n_51680_65240 Rseg
X2611 n_51680_65240 n_51680_68040 Rseg
X2612 n_51680_68040 n_51680_70840 Rseg
X2613 n_51680_70840 n_51680_73640 Rseg
X2614 n_51680_73640 n_51680_76440 Rseg
X2615 n_51680_76440 n_51680_79240 Rseg
X2616 n_51680_79240 n_51680_82040 Rseg
X2617 n_51680_82040 n_51680_84840 Rseg
X2618 n_51680_84840 n_51680_87640 Rseg
X2619 n_52060_40040 n_52060_42840 Rseg
X2620 n_52060_42840 n_52060_45640 Rseg
X2621 n_52060_45640 n_52060_48440 Rseg
X2622 n_52060_48440 n_52060_51240 Rseg
X2623 n_52060_51240 n_52060_54040 Rseg
X2624 n_52060_54040 n_52060_56840 Rseg
X2625 n_52060_56840 n_52060_59640 Rseg
X2626 n_52060_59640 n_52060_62440 Rseg
X2627 n_52060_62440 n_52060_65240 Rseg
X2628 n_52060_65240 n_52060_68040 Rseg
X2629 n_52060_68040 n_52060_70840 Rseg
X2630 n_52060_70840 n_52060_73640 Rseg
X2631 n_52060_73640 n_52060_76440 Rseg
X2632 n_52060_76440 n_52060_79240 Rseg
X2633 n_52060_79240 n_52060_82040 Rseg
X2634 n_52060_82040 n_52060_84840 Rseg
X2635 n_52060_84840 n_52060_87640 Rseg
X2636 n_52440_40040 n_52440_42840 Rseg
X2637 n_52440_42840 n_52440_45640 Rseg
X2638 n_52440_45640 n_52440_48440 Rseg
X2639 n_52440_48440 n_52440_51240 Rseg
X2640 n_52440_51240 n_52440_54040 Rseg
X2641 n_52440_54040 n_52440_56840 Rseg
X2642 n_52440_56840 n_52440_59640 Rseg
X2643 n_52440_59640 n_52440_62440 Rseg
X2644 n_52440_62440 n_52440_65240 Rseg
X2645 n_52440_65240 n_52440_68040 Rseg
X2646 n_52440_68040 n_52440_70840 Rseg
X2647 n_52440_70840 n_52440_73640 Rseg
X2648 n_52440_73640 n_52440_76440 Rseg
X2649 n_52440_76440 n_52440_79240 Rseg
X2650 n_52440_79240 n_52440_82040 Rseg
X2651 n_52440_82040 n_52440_84840 Rseg
X2652 n_52440_84840 n_52440_87640 Rseg
X2653 n_52820_40040 n_52820_42840 Rseg
X2654 n_52820_42840 n_52820_45640 Rseg
X2655 n_52820_45640 n_52820_48440 Rseg
X2656 n_52820_48440 n_52820_51240 Rseg
X2657 n_52820_51240 n_52820_54040 Rseg
X2658 n_52820_54040 n_52820_56840 Rseg
X2659 n_52820_56840 n_52820_59640 Rseg
X2660 n_52820_59640 n_52820_62440 Rseg
X2661 n_52820_62440 n_52820_65240 Rseg
X2662 n_52820_65240 n_52820_68040 Rseg
X2663 n_52820_68040 n_52820_70840 Rseg
X2664 n_52820_70840 n_52820_73640 Rseg
X2665 n_52820_73640 n_52820_76440 Rseg
X2666 n_52820_76440 n_52820_79240 Rseg
X2667 n_52820_79240 n_52820_82040 Rseg
X2668 n_52820_82040 n_52820_84840 Rseg
X2669 n_52820_84840 n_52820_87640 Rseg
X2670 n_53200_40040 n_53200_42840 Rseg
X2671 n_53200_42840 n_53200_45640 Rseg
X2672 n_53200_45640 n_53200_48440 Rseg
X2673 n_53200_48440 n_53200_51240 Rseg
X2674 n_53200_51240 n_53200_54040 Rseg
X2675 n_53200_54040 n_53200_56840 Rseg
X2676 n_53200_56840 n_53200_59640 Rseg
X2677 n_53200_59640 n_53200_62440 Rseg
X2678 n_53200_62440 n_53200_65240 Rseg
X2679 n_53200_65240 n_53200_68040 Rseg
X2680 n_53200_68040 n_53200_70840 Rseg
X2681 n_53200_70840 n_53200_73640 Rseg
X2682 n_53200_73640 n_53200_76440 Rseg
X2683 n_53200_76440 n_53200_79240 Rseg
X2684 n_53200_79240 n_53200_82040 Rseg
X2685 n_53200_82040 n_53200_84840 Rseg
X2686 n_53200_84840 n_53200_87640 Rseg
X2687 n_53580_40040 n_53580_42840 Rseg
X2688 n_53580_42840 n_53580_45640 Rseg
X2689 n_53580_45640 n_53580_48440 Rseg
X2690 n_53580_48440 n_53580_51240 Rseg
X2691 n_53580_51240 n_53580_54040 Rseg
X2692 n_53580_54040 n_53580_56840 Rseg
X2693 n_53580_56840 n_53580_59640 Rseg
X2694 n_53580_59640 n_53580_62440 Rseg
X2695 n_53580_62440 n_53580_65240 Rseg
X2696 n_53580_65240 n_53580_68040 Rseg
X2697 n_53580_68040 n_53580_70840 Rseg
X2698 n_53580_70840 n_53580_73640 Rseg
X2699 n_53580_73640 n_53580_76440 Rseg
X2700 n_53580_76440 n_53580_79240 Rseg
X2701 n_53580_79240 n_53580_82040 Rseg
X2702 n_53580_82040 n_53580_84840 Rseg
X2703 n_53580_84840 n_53580_87640 Rseg
X2704 n_53960_40040 n_53960_42840 Rseg
X2705 n_53960_42840 n_53960_45640 Rseg
X2706 n_53960_45640 n_53960_48440 Rseg
X2707 n_53960_48440 n_53960_51240 Rseg
X2708 n_53960_51240 n_53960_54040 Rseg
X2709 n_53960_54040 n_53960_56840 Rseg
X2710 n_53960_56840 n_53960_59640 Rseg
X2711 n_53960_59640 n_53960_62440 Rseg
X2712 n_53960_62440 n_53960_65240 Rseg
X2713 n_53960_65240 n_53960_68040 Rseg
X2714 n_53960_68040 n_53960_70840 Rseg
X2715 n_53960_70840 n_53960_73640 Rseg
X2716 n_53960_73640 n_53960_76440 Rseg
X2717 n_53960_76440 n_53960_79240 Rseg
X2718 n_53960_79240 n_53960_82040 Rseg
X2719 n_53960_82040 n_53960_84840 Rseg
X2720 n_53960_84840 n_53960_87640 Rseg
X2721 n_54340_40040 n_54340_42840 Rseg
X2722 n_54340_42840 n_54340_45640 Rseg
X2723 n_54340_45640 n_54340_48440 Rseg
X2724 n_54340_48440 n_54340_51240 Rseg
X2725 n_54340_51240 n_54340_54040 Rseg
X2726 n_54340_54040 n_54340_56840 Rseg
X2727 n_54340_56840 n_54340_59640 Rseg
X2728 n_54340_59640 n_54340_62440 Rseg
X2729 n_54340_62440 n_54340_65240 Rseg
X2730 n_54340_65240 n_54340_68040 Rseg
X2731 n_54340_68040 n_54340_70840 Rseg
X2732 n_54340_70840 n_54340_73640 Rseg
X2733 n_54340_73640 n_54340_76440 Rseg
X2734 n_54340_76440 n_54340_79240 Rseg
X2735 n_54340_79240 n_54340_82040 Rseg
X2736 n_54340_82040 n_54340_84840 Rseg
X2737 n_54340_84840 n_54340_87640 Rseg
X2738 n_54720_40040 n_54720_42840 Rseg
X2739 n_54720_42840 n_54720_45640 Rseg
X2740 n_54720_45640 n_54720_48440 Rseg
X2741 n_54720_48440 n_54720_51240 Rseg
X2742 n_54720_51240 n_54720_54040 Rseg
X2743 n_54720_54040 n_54720_56840 Rseg
X2744 n_54720_56840 n_54720_59640 Rseg
X2745 n_54720_59640 n_54720_62440 Rseg
X2746 n_54720_62440 n_54720_65240 Rseg
X2747 n_54720_65240 n_54720_68040 Rseg
X2748 n_54720_68040 n_54720_70840 Rseg
X2749 n_54720_70840 n_54720_73640 Rseg
X2750 n_54720_73640 n_54720_76440 Rseg
X2751 n_54720_76440 n_54720_79240 Rseg
X2752 n_54720_79240 n_54720_82040 Rseg
X2753 n_54720_82040 n_54720_84840 Rseg
X2754 n_54720_84840 n_54720_87640 Rseg
X2755 n_55100_40040 n_55100_42840 Rseg
X2756 n_55100_42840 n_55100_45640 Rseg
X2757 n_55100_45640 n_55100_48440 Rseg
X2758 n_55100_48440 n_55100_51240 Rseg
X2759 n_55100_51240 n_55100_54040 Rseg
X2760 n_55100_54040 n_55100_56840 Rseg
X2761 n_55100_56840 n_55100_59640 Rseg
X2762 n_55100_59640 n_55100_62440 Rseg
X2763 n_55100_62440 n_55100_65240 Rseg
X2764 n_55100_65240 n_55100_68040 Rseg
X2765 n_55100_68040 n_55100_70840 Rseg
X2766 n_55100_70840 n_55100_73640 Rseg
X2767 n_55100_73640 n_55100_76440 Rseg
X2768 n_55100_76440 n_55100_79240 Rseg
X2769 n_55100_79240 n_55100_82040 Rseg
X2770 n_55100_82040 n_55100_84840 Rseg
X2771 n_55100_84840 n_55100_87640 Rseg
X2772 n_55480_40040 n_55480_42840 Rseg
X2773 n_55480_42840 n_55480_45640 Rseg
X2774 n_55480_45640 n_55480_48440 Rseg
X2775 n_55480_48440 n_55480_51240 Rseg
X2776 n_55480_51240 n_55480_54040 Rseg
X2777 n_55480_54040 n_55480_56840 Rseg
X2778 n_55480_56840 n_55480_59640 Rseg
X2779 n_55480_59640 n_55480_62440 Rseg
X2780 n_55480_62440 n_55480_65240 Rseg
X2781 n_55480_65240 n_55480_68040 Rseg
X2782 n_55480_68040 n_55480_70840 Rseg
X2783 n_55480_70840 n_55480_73640 Rseg
X2784 n_55480_73640 n_55480_76440 Rseg
X2785 n_55480_76440 n_55480_79240 Rseg
X2786 n_55480_79240 n_55480_82040 Rseg
X2787 n_55480_82040 n_55480_84840 Rseg
X2788 n_55480_84840 n_55480_87640 Rseg
X2789 n_55860_40040 n_55860_42840 Rseg
X2790 n_55860_42840 n_55860_45640 Rseg
X2791 n_55860_45640 n_55860_48440 Rseg
X2792 n_55860_48440 n_55860_51240 Rseg
X2793 n_55860_51240 n_55860_54040 Rseg
X2794 n_55860_54040 n_55860_56840 Rseg
X2795 n_55860_56840 n_55860_59640 Rseg
X2796 n_55860_59640 n_55860_62440 Rseg
X2797 n_55860_62440 n_55860_65240 Rseg
X2798 n_55860_65240 n_55860_68040 Rseg
X2799 n_55860_68040 n_55860_70840 Rseg
X2800 n_55860_70840 n_55860_73640 Rseg
X2801 n_55860_73640 n_55860_76440 Rseg
X2802 n_55860_76440 n_55860_79240 Rseg
X2803 n_55860_79240 n_55860_82040 Rseg
X2804 n_55860_82040 n_55860_84840 Rseg
X2805 n_55860_84840 n_55860_87640 Rseg
X2806 n_56240_40040 n_56240_42840 Rseg
X2807 n_56240_42840 n_56240_45640 Rseg
X2808 n_56240_45640 n_56240_48440 Rseg
X2809 n_56240_48440 n_56240_51240 Rseg
X2810 n_56240_51240 n_56240_54040 Rseg
X2811 n_56240_54040 n_56240_56840 Rseg
X2812 n_56240_56840 n_56240_59640 Rseg
X2813 n_56240_59640 n_56240_62440 Rseg
X2814 n_56240_62440 n_56240_65240 Rseg
X2815 n_56240_65240 n_56240_68040 Rseg
X2816 n_56240_68040 n_56240_70840 Rseg
X2817 n_56240_70840 n_56240_73640 Rseg
X2818 n_56240_73640 n_56240_76440 Rseg
X2819 n_56240_76440 n_56240_79240 Rseg
X2820 n_56240_79240 n_56240_82040 Rseg
X2821 n_56240_82040 n_56240_84840 Rseg
X2822 n_56240_84840 n_56240_87640 Rseg
X2823 n_56620_40040 n_56620_42840 Rseg
X2824 n_56620_42840 n_56620_45640 Rseg
X2825 n_56620_45640 n_56620_48440 Rseg
X2826 n_56620_48440 n_56620_51240 Rseg
X2827 n_56620_51240 n_56620_54040 Rseg
X2828 n_56620_54040 n_56620_56840 Rseg
X2829 n_56620_56840 n_56620_59640 Rseg
X2830 n_56620_59640 n_56620_62440 Rseg
X2831 n_56620_62440 n_56620_65240 Rseg
X2832 n_56620_65240 n_56620_68040 Rseg
X2833 n_56620_68040 n_56620_70840 Rseg
X2834 n_56620_70840 n_56620_73640 Rseg
X2835 n_56620_73640 n_56620_76440 Rseg
X2836 n_56620_76440 n_56620_79240 Rseg
X2837 n_56620_79240 n_56620_82040 Rseg
X2838 n_56620_82040 n_56620_84840 Rseg
X2839 n_56620_84840 n_56620_87640 Rseg
X2840 n_57000_40040 n_57000_42840 Rseg
X2841 n_57000_42840 n_57000_45640 Rseg
X2842 n_57000_45640 n_57000_48440 Rseg
X2843 n_57000_48440 n_57000_51240 Rseg
X2844 n_57000_51240 n_57000_54040 Rseg
X2845 n_57000_54040 n_57000_56840 Rseg
X2846 n_57000_56840 n_57000_59640 Rseg
X2847 n_57000_59640 n_57000_62440 Rseg
X2848 n_57000_62440 n_57000_65240 Rseg
X2849 n_57000_65240 n_57000_68040 Rseg
X2850 n_57000_68040 n_57000_70840 Rseg
X2851 n_57000_70840 n_57000_73640 Rseg
X2852 n_57000_73640 n_57000_76440 Rseg
X2853 n_57000_76440 n_57000_79240 Rseg
X2854 n_57000_79240 n_57000_82040 Rseg
X2855 n_57000_82040 n_57000_84840 Rseg
X2856 n_57000_84840 n_57000_87640 Rseg
X2857 n_57380_40040 n_57380_42840 Rseg
X2858 n_57380_42840 n_57380_45640 Rseg
X2859 n_57380_45640 n_57380_48440 Rseg
X2860 n_57380_48440 n_57380_51240 Rseg
X2861 n_57380_51240 n_57380_54040 Rseg
X2862 n_57380_54040 n_57380_56840 Rseg
X2863 n_57380_56840 n_57380_59640 Rseg
X2864 n_57380_59640 n_57380_62440 Rseg
X2865 n_57380_62440 n_57380_65240 Rseg
X2866 n_57380_65240 n_57380_68040 Rseg
X2867 n_57380_68040 n_57380_70840 Rseg
X2868 n_57380_70840 n_57380_73640 Rseg
X2869 n_57380_73640 n_57380_76440 Rseg
X2870 n_57380_76440 n_57380_79240 Rseg
X2871 n_57380_79240 n_57380_82040 Rseg
X2872 n_57380_82040 n_57380_84840 Rseg
X2873 n_57380_84840 n_57380_87640 Rseg
X2874 n_57760_40040 n_57760_42840 Rseg
X2875 n_57760_42840 n_57760_45640 Rseg
X2876 n_57760_45640 n_57760_48440 Rseg
X2877 n_57760_48440 n_57760_51240 Rseg
X2878 n_57760_51240 n_57760_54040 Rseg
X2879 n_57760_54040 n_57760_56840 Rseg
X2880 n_57760_56840 n_57760_59640 Rseg
X2881 n_57760_59640 n_57760_62440 Rseg
X2882 n_57760_62440 n_57760_65240 Rseg
X2883 n_57760_65240 n_57760_68040 Rseg
X2884 n_57760_68040 n_57760_70840 Rseg
X2885 n_57760_70840 n_57760_73640 Rseg
X2886 n_57760_73640 n_57760_76440 Rseg
X2887 n_57760_76440 n_57760_79240 Rseg
X2888 n_57760_79240 n_57760_82040 Rseg
X2889 n_57760_82040 n_57760_84840 Rseg
X2890 n_57760_84840 n_57760_87640 Rseg
X2891 n_58140_40040 n_58140_42840 Rseg
X2892 n_58140_42840 n_58140_45640 Rseg
X2893 n_58140_45640 n_58140_48440 Rseg
X2894 n_58140_48440 n_58140_51240 Rseg
X2895 n_58140_51240 n_58140_54040 Rseg
X2896 n_58140_54040 n_58140_56840 Rseg
X2897 n_58140_56840 n_58140_59640 Rseg
X2898 n_58140_59640 n_58140_62440 Rseg
X2899 n_58140_62440 n_58140_65240 Rseg
X2900 n_58140_65240 n_58140_68040 Rseg
X2901 n_58140_68040 n_58140_70840 Rseg
X2902 n_58140_70840 n_58140_73640 Rseg
X2903 n_58140_73640 n_58140_76440 Rseg
X2904 n_58140_76440 n_58140_79240 Rseg
X2905 n_58140_79240 n_58140_82040 Rseg
X2906 n_58140_82040 n_58140_84840 Rseg
X2907 n_58140_84840 n_58140_87640 Rseg
X2908 n_58520_40040 n_58520_42840 Rseg
X2909 n_58520_42840 n_58520_45640 Rseg
X2910 n_58520_45640 n_58520_48440 Rseg
X2911 n_58520_48440 n_58520_51240 Rseg
X2912 n_58520_51240 n_58520_54040 Rseg
X2913 n_58520_54040 n_58520_56840 Rseg
X2914 n_58520_56840 n_58520_59640 Rseg
X2915 n_58520_59640 n_58520_62440 Rseg
X2916 n_58520_62440 n_58520_65240 Rseg
X2917 n_58520_65240 n_58520_68040 Rseg
X2918 n_58520_68040 n_58520_70840 Rseg
X2919 n_58520_70840 n_58520_73640 Rseg
X2920 n_58520_73640 n_58520_76440 Rseg
X2921 n_58520_76440 n_58520_79240 Rseg
X2922 n_58520_79240 n_58520_82040 Rseg
X2923 n_58520_82040 n_58520_84840 Rseg
X2924 n_58520_84840 n_58520_87640 Rseg
X2925 n_58900_40040 n_58900_42840 Rseg
X2926 n_58900_42840 n_58900_45640 Rseg
X2927 n_58900_45640 n_58900_48440 Rseg
X2928 n_58900_48440 n_58900_51240 Rseg
X2929 n_58900_51240 n_58900_54040 Rseg
X2930 n_58900_54040 n_58900_56840 Rseg
X2931 n_58900_56840 n_58900_59640 Rseg
X2932 n_58900_59640 n_58900_62440 Rseg
X2933 n_58900_62440 n_58900_65240 Rseg
X2934 n_58900_65240 n_58900_68040 Rseg
X2935 n_58900_68040 n_58900_70840 Rseg
X2936 n_58900_70840 n_58900_73640 Rseg
X2937 n_58900_73640 n_58900_76440 Rseg
X2938 n_58900_76440 n_58900_79240 Rseg
X2939 n_58900_79240 n_58900_82040 Rseg
X2940 n_58900_82040 n_58900_84840 Rseg
X2941 n_58900_84840 n_58900_87640 Rseg
X2942 n_59280_40040 n_59280_42840 Rseg
X2943 n_59280_42840 n_59280_45640 Rseg
X2944 n_59280_45640 n_59280_48440 Rseg
X2945 n_59280_48440 n_59280_51240 Rseg
X2946 n_59280_51240 n_59280_54040 Rseg
X2947 n_59280_54040 n_59280_56840 Rseg
X2948 n_59280_56840 n_59280_59640 Rseg
X2949 n_59280_59640 n_59280_62440 Rseg
X2950 n_59280_62440 n_59280_65240 Rseg
X2951 n_59280_65240 n_59280_68040 Rseg
X2952 n_59280_68040 n_59280_70840 Rseg
X2953 n_59280_70840 n_59280_73640 Rseg
X2954 n_59280_73640 n_59280_76440 Rseg
X2955 n_59280_76440 n_59280_79240 Rseg
X2956 n_59280_79240 n_59280_82040 Rseg
X2957 n_59280_82040 n_59280_84840 Rseg
X2958 n_59280_84840 n_59280_87640 Rseg
X2959 n_59660_40040 n_59660_42840 Rseg
X2960 n_59660_42840 n_59660_45640 Rseg
X2961 n_59660_45640 n_59660_48440 Rseg
X2962 n_59660_48440 n_59660_51240 Rseg
X2963 n_59660_51240 n_59660_54040 Rseg
X2964 n_59660_54040 n_59660_56840 Rseg
X2965 n_59660_56840 n_59660_59640 Rseg
X2966 n_59660_59640 n_59660_62440 Rseg
X2967 n_59660_62440 n_59660_65240 Rseg
X2968 n_59660_65240 n_59660_68040 Rseg
X2969 n_59660_68040 n_59660_70840 Rseg
X2970 n_59660_70840 n_59660_73640 Rseg
X2971 n_59660_73640 n_59660_76440 Rseg
X2972 n_59660_76440 n_59660_79240 Rseg
X2973 n_59660_79240 n_59660_82040 Rseg
X2974 n_59660_82040 n_59660_84840 Rseg
X2975 n_59660_84840 n_59660_87640 Rseg
X2976 n_60040_40040 n_60040_42840 Rseg
X2977 n_60040_42840 n_60040_45640 Rseg
X2978 n_60040_45640 n_60040_48440 Rseg
X2979 n_60040_48440 n_60040_51240 Rseg
X2980 n_60040_51240 n_60040_54040 Rseg
X2981 n_60040_54040 n_60040_56840 Rseg
X2982 n_60040_56840 n_60040_59640 Rseg
X2983 n_60040_59640 n_60040_62440 Rseg
X2984 n_60040_62440 n_60040_65240 Rseg
X2985 n_60040_65240 n_60040_68040 Rseg
X2986 n_60040_68040 n_60040_70840 Rseg
X2987 n_60040_70840 n_60040_73640 Rseg
X2988 n_60040_73640 n_60040_76440 Rseg
X2989 n_60040_76440 n_60040_79240 Rseg
X2990 n_60040_79240 n_60040_82040 Rseg
X2991 n_60040_82040 n_60040_84840 Rseg
X2992 n_60040_84840 n_60040_87640 Rseg
X2993 n_60420_40040 n_60420_42840 Rseg
X2994 n_60420_42840 n_60420_45640 Rseg
X2995 n_60420_45640 n_60420_48440 Rseg
X2996 n_60420_48440 n_60420_51240 Rseg
X2997 n_60420_51240 n_60420_54040 Rseg
X2998 n_60420_54040 n_60420_56840 Rseg
X2999 n_60420_56840 n_60420_59640 Rseg
X3000 n_60420_59640 n_60420_62440 Rseg
X3001 n_60420_62440 n_60420_65240 Rseg
X3002 n_60420_65240 n_60420_68040 Rseg
X3003 n_60420_68040 n_60420_70840 Rseg
X3004 n_60420_70840 n_60420_73640 Rseg
X3005 n_60420_73640 n_60420_76440 Rseg
X3006 n_60420_76440 n_60420_79240 Rseg
X3007 n_60420_79240 n_60420_82040 Rseg
X3008 n_60420_82040 n_60420_84840 Rseg
X3009 n_60420_84840 n_60420_87640 Rseg
X3010 n_60800_40040 n_60800_42840 Rseg
X3011 n_60800_42840 n_60800_45640 Rseg
X3012 n_60800_45640 n_60800_48440 Rseg
X3013 n_60800_48440 n_60800_51240 Rseg
X3014 n_60800_51240 n_60800_54040 Rseg
X3015 n_60800_54040 n_60800_56840 Rseg
X3016 n_60800_56840 n_60800_59640 Rseg
X3017 n_60800_59640 n_60800_62440 Rseg
X3018 n_60800_62440 n_60800_65240 Rseg
X3019 n_60800_65240 n_60800_68040 Rseg
X3020 n_60800_68040 n_60800_70840 Rseg
X3021 n_60800_70840 n_60800_73640 Rseg
X3022 n_60800_73640 n_60800_76440 Rseg
X3023 n_60800_76440 n_60800_79240 Rseg
X3024 n_60800_79240 n_60800_82040 Rseg
X3025 n_60800_82040 n_60800_84840 Rseg
X3026 n_60800_84840 n_60800_87640 Rseg
X3027 n_61180_40040 n_61180_42840 Rseg
X3028 n_61180_42840 n_61180_45640 Rseg
X3029 n_61180_45640 n_61180_48440 Rseg
X3030 n_61180_48440 n_61180_51240 Rseg
X3031 n_61180_51240 n_61180_54040 Rseg
X3032 n_61180_54040 n_61180_56840 Rseg
X3033 n_61180_56840 n_61180_59640 Rseg
X3034 n_61180_59640 n_61180_62440 Rseg
X3035 n_61180_62440 n_61180_65240 Rseg
X3036 n_61180_65240 n_61180_68040 Rseg
X3037 n_61180_68040 n_61180_70840 Rseg
X3038 n_61180_70840 n_61180_73640 Rseg
X3039 n_61180_73640 n_61180_76440 Rseg
X3040 n_61180_76440 n_61180_79240 Rseg
X3041 n_61180_79240 n_61180_82040 Rseg
X3042 n_61180_82040 n_61180_84840 Rseg
X3043 n_61180_84840 n_61180_87640 Rseg
X3044 n_61560_40040 n_61560_42840 Rseg
X3045 n_61560_42840 n_61560_45640 Rseg
X3046 n_61560_45640 n_61560_48440 Rseg
X3047 n_61560_48440 n_61560_51240 Rseg
X3048 n_61560_51240 n_61560_54040 Rseg
X3049 n_61560_54040 n_61560_56840 Rseg
X3050 n_61560_56840 n_61560_59640 Rseg
X3051 n_61560_59640 n_61560_62440 Rseg
X3052 n_61560_62440 n_61560_65240 Rseg
X3053 n_61560_65240 n_61560_68040 Rseg
X3054 n_61560_68040 n_61560_70840 Rseg
X3055 n_61560_70840 n_61560_73640 Rseg
X3056 n_61560_73640 n_61560_76440 Rseg
X3057 n_61560_76440 n_61560_79240 Rseg
X3058 n_61560_79240 n_61560_82040 Rseg
X3059 n_61560_82040 n_61560_84840 Rseg
X3060 n_61560_84840 n_61560_87640 Rseg
X3061 n_61940_40040 n_61940_42840 Rseg
X3062 n_61940_42840 n_61940_45640 Rseg
X3063 n_61940_45640 n_61940_48440 Rseg
X3064 n_61940_48440 n_61940_51240 Rseg
X3065 n_61940_51240 n_61940_54040 Rseg
X3066 n_61940_54040 n_61940_56840 Rseg
X3067 n_61940_56840 n_61940_59640 Rseg
X3068 n_61940_59640 n_61940_62440 Rseg
X3069 n_61940_62440 n_61940_65240 Rseg
X3070 n_61940_65240 n_61940_68040 Rseg
X3071 n_61940_68040 n_61940_70840 Rseg
X3072 n_61940_70840 n_61940_73640 Rseg
X3073 n_61940_73640 n_61940_76440 Rseg
X3074 n_61940_76440 n_61940_79240 Rseg
X3075 n_61940_79240 n_61940_82040 Rseg
X3076 n_61940_82040 n_61940_84840 Rseg
X3077 n_61940_84840 n_61940_87640 Rseg
X3078 n_62320_40040 n_62320_42840 Rseg
X3079 n_62320_42840 n_62320_45640 Rseg
X3080 n_62320_45640 n_62320_48440 Rseg
X3081 n_62320_48440 n_62320_51240 Rseg
X3082 n_62320_51240 n_62320_54040 Rseg
X3083 n_62320_54040 n_62320_56840 Rseg
X3084 n_62320_56840 n_62320_59640 Rseg
X3085 n_62320_59640 n_62320_62440 Rseg
X3086 n_62320_62440 n_62320_65240 Rseg
X3087 n_62320_65240 n_62320_68040 Rseg
X3088 n_62320_68040 n_62320_70840 Rseg
X3089 n_62320_70840 n_62320_73640 Rseg
X3090 n_62320_73640 n_62320_76440 Rseg
X3091 n_62320_76440 n_62320_79240 Rseg
X3092 n_62320_79240 n_62320_82040 Rseg
X3093 n_62320_82040 n_62320_84840 Rseg
X3094 n_62320_84840 n_62320_87640 Rseg
X3095 n_63080_40040 n_63080_42840 Rseg
X3096 n_63080_42840 n_63080_45640 Rseg
X3097 n_63080_45640 n_63080_48440 Rseg
X3098 n_63080_48440 n_63080_51240 Rseg
X3099 n_63080_51240 n_63080_54040 Rseg
X3100 n_63080_54040 n_63080_56840 Rseg
X3101 n_63080_56840 n_63080_59640 Rseg
X3102 n_63080_59640 n_63080_62440 Rseg
X3103 n_63080_62440 n_63080_65240 Rseg
X3104 n_63080_65240 n_63080_68040 Rseg
X3105 n_63080_68040 n_63080_70840 Rseg
X3106 n_63080_70840 n_63080_73640 Rseg
X3107 n_63080_73640 n_63080_76440 Rseg
X3108 n_63080_76440 n_63080_79240 Rseg
X3109 n_63080_79240 n_63080_82040 Rseg
X3110 n_63080_82040 n_63080_84840 Rseg
X3111 n_63080_84840 n_63080_87640 Rseg
X3112 n_63460_40040 n_63460_42840 Rseg
X3113 n_63460_42840 n_63460_45640 Rseg
X3114 n_63460_45640 n_63460_48440 Rseg
X3115 n_63460_48440 n_63460_51240 Rseg
X3116 n_63460_51240 n_63460_54040 Rseg
X3117 n_63460_54040 n_63460_56840 Rseg
X3118 n_63460_56840 n_63460_59640 Rseg
X3119 n_63460_59640 n_63460_62440 Rseg
X3120 n_63460_62440 n_63460_65240 Rseg
X3121 n_63460_65240 n_63460_68040 Rseg
X3122 n_63460_68040 n_63460_70840 Rseg
X3123 n_63460_70840 n_63460_73640 Rseg
X3124 n_63460_73640 n_63460_76440 Rseg
X3125 n_63460_76440 n_63460_79240 Rseg
X3126 n_63460_79240 n_63460_82040 Rseg
X3127 n_63460_82040 n_63460_84840 Rseg
X3128 n_63460_84840 n_63460_87640 Rseg
X3129 n_63840_40040 n_63840_42840 Rseg
X3130 n_63840_42840 n_63840_45640 Rseg
X3131 n_63840_45640 n_63840_48440 Rseg
X3132 n_63840_48440 n_63840_51240 Rseg
X3133 n_63840_51240 n_63840_54040 Rseg
X3134 n_63840_54040 n_63840_56840 Rseg
X3135 n_63840_56840 n_63840_59640 Rseg
X3136 n_63840_59640 n_63840_62440 Rseg
X3137 n_63840_62440 n_63840_65240 Rseg
X3138 n_63840_65240 n_63840_68040 Rseg
X3139 n_63840_68040 n_63840_70840 Rseg
X3140 n_63840_70840 n_63840_73640 Rseg
X3141 n_63840_73640 n_63840_76440 Rseg
X3142 n_63840_76440 n_63840_79240 Rseg
X3143 n_63840_79240 n_63840_82040 Rseg
X3144 n_63840_82040 n_63840_84840 Rseg
X3145 n_63840_84840 n_63840_87640 Rseg
X3146 n_64220_40040 n_64220_42840 Rseg
X3147 n_64220_42840 n_64220_45640 Rseg
X3148 n_64220_45640 n_64220_48440 Rseg
X3149 n_64220_48440 n_64220_51240 Rseg
X3150 n_64220_51240 n_64220_54040 Rseg
X3151 n_64220_54040 n_64220_56840 Rseg
X3152 n_64220_56840 n_64220_59640 Rseg
X3153 n_64220_59640 n_64220_62440 Rseg
X3154 n_64220_62440 n_64220_65240 Rseg
X3155 n_64220_65240 n_64220_68040 Rseg
X3156 n_64220_68040 n_64220_70840 Rseg
X3157 n_64220_70840 n_64220_73640 Rseg
X3158 n_64220_73640 n_64220_76440 Rseg
X3159 n_64220_76440 n_64220_79240 Rseg
X3160 n_64220_79240 n_64220_82040 Rseg
X3161 n_64220_82040 n_64220_84840 Rseg
X3162 n_64220_84840 n_64220_87640 Rseg
X3163 n_64600_40040 n_64600_42840 Rseg
X3164 n_64600_42840 n_64600_45640 Rseg
X3165 n_64600_45640 n_64600_48440 Rseg
X3166 n_64600_48440 n_64600_51240 Rseg
X3167 n_64600_51240 n_64600_54040 Rseg
X3168 n_64600_54040 n_64600_56840 Rseg
X3169 n_64600_56840 n_64600_59640 Rseg
X3170 n_64600_59640 n_64600_62440 Rseg
X3171 n_64600_62440 n_64600_65240 Rseg
X3172 n_64600_65240 n_64600_68040 Rseg
X3173 n_64600_68040 n_64600_70840 Rseg
X3174 n_64600_70840 n_64600_73640 Rseg
X3175 n_64600_73640 n_64600_76440 Rseg
X3176 n_64600_76440 n_64600_79240 Rseg
X3177 n_64600_79240 n_64600_82040 Rseg
X3178 n_64600_82040 n_64600_84840 Rseg
X3179 n_64600_84840 n_64600_87640 Rseg
X3180 n_64980_40040 n_64980_42840 Rseg
X3181 n_64980_42840 n_64980_45640 Rseg
X3182 n_64980_45640 n_64980_48440 Rseg
X3183 n_64980_48440 n_64980_51240 Rseg
X3184 n_64980_51240 n_64980_54040 Rseg
X3185 n_64980_54040 n_64980_56840 Rseg
X3186 n_64980_56840 n_64980_59640 Rseg
X3187 n_64980_59640 n_64980_62440 Rseg
X3188 n_64980_62440 n_64980_65240 Rseg
X3189 n_64980_65240 n_64980_68040 Rseg
X3190 n_64980_68040 n_64980_70840 Rseg
X3191 n_64980_70840 n_64980_73640 Rseg
X3192 n_64980_73640 n_64980_76440 Rseg
X3193 n_64980_76440 n_64980_79240 Rseg
X3194 n_64980_79240 n_64980_82040 Rseg
X3195 n_64980_82040 n_64980_84840 Rseg
X3196 n_64980_84840 n_64980_87640 Rseg
X3197 n_65360_40040 n_65360_42840 Rseg
X3198 n_65360_42840 n_65360_45640 Rseg
X3199 n_65360_45640 n_65360_48440 Rseg
X3200 n_65360_48440 n_65360_51240 Rseg
X3201 n_65360_51240 n_65360_54040 Rseg
X3202 n_65360_54040 n_65360_56840 Rseg
X3203 n_65360_56840 n_65360_59640 Rseg
X3204 n_65360_59640 n_65360_62440 Rseg
X3205 n_65360_62440 n_65360_65240 Rseg
X3206 n_65360_65240 n_65360_68040 Rseg
X3207 n_65360_68040 n_65360_70840 Rseg
X3208 n_65360_70840 n_65360_73640 Rseg
X3209 n_65360_73640 n_65360_76440 Rseg
X3210 n_65360_76440 n_65360_79240 Rseg
X3211 n_65360_79240 n_65360_82040 Rseg
X3212 n_65360_82040 n_65360_84840 Rseg
X3213 n_65360_84840 n_65360_87640 Rseg
X3214 n_65740_40040 n_65740_42840 Rseg
X3215 n_65740_42840 n_65740_45640 Rseg
X3216 n_65740_45640 n_65740_48440 Rseg
X3217 n_65740_48440 n_65740_51240 Rseg
X3218 n_65740_51240 n_65740_54040 Rseg
X3219 n_65740_54040 n_65740_56840 Rseg
X3220 n_65740_56840 n_65740_59640 Rseg
X3221 n_65740_59640 n_65740_62440 Rseg
X3222 n_65740_62440 n_65740_65240 Rseg
X3223 n_65740_65240 n_65740_68040 Rseg
X3224 n_65740_68040 n_65740_70840 Rseg
X3225 n_65740_70840 n_65740_73640 Rseg
X3226 n_65740_73640 n_65740_76440 Rseg
X3227 n_65740_76440 n_65740_79240 Rseg
X3228 n_65740_79240 n_65740_82040 Rseg
X3229 n_65740_82040 n_65740_84840 Rseg
X3230 n_65740_84840 n_65740_87640 Rseg
X3231 n_66120_40040 n_66120_42840 Rseg
X3232 n_66120_42840 n_66120_45640 Rseg
X3233 n_66120_45640 n_66120_48440 Rseg
X3234 n_66120_48440 n_66120_51240 Rseg
X3235 n_66120_51240 n_66120_54040 Rseg
X3236 n_66120_54040 n_66120_56840 Rseg
X3237 n_66120_56840 n_66120_59640 Rseg
X3238 n_66120_59640 n_66120_62440 Rseg
X3239 n_66120_62440 n_66120_65240 Rseg
X3240 n_66120_65240 n_66120_68040 Rseg
X3241 n_66120_68040 n_66120_70840 Rseg
X3242 n_66120_70840 n_66120_73640 Rseg
X3243 n_66120_73640 n_66120_76440 Rseg
X3244 n_66120_76440 n_66120_79240 Rseg
X3245 n_66120_79240 n_66120_82040 Rseg
X3246 n_66120_82040 n_66120_84840 Rseg
X3247 n_66120_84840 n_66120_87640 Rseg
X3248 n_66880_40040 n_66880_42840 Rseg
X3249 n_66880_42840 n_66880_45640 Rseg
X3250 n_66880_45640 n_66880_48440 Rseg
X3251 n_66880_48440 n_66880_51240 Rseg
X3252 n_66880_51240 n_66880_54040 Rseg
X3253 n_66880_54040 n_66880_56840 Rseg
X3254 n_66880_56840 n_66880_59640 Rseg
X3255 n_66880_59640 n_66880_62440 Rseg
X3256 n_66880_62440 n_66880_65240 Rseg
X3257 n_66880_65240 n_66880_68040 Rseg
X3258 n_66880_68040 n_66880_70840 Rseg
X3259 n_66880_70840 n_66880_73640 Rseg
X3260 n_66880_73640 n_66880_76440 Rseg
X3261 n_66880_76440 n_66880_79240 Rseg
X3262 n_66880_79240 n_66880_82040 Rseg
X3263 n_66880_82040 n_66880_84840 Rseg
X3264 n_66880_84840 n_66880_87640 Rseg
X3265 n_67260_40040 n_67260_42840 Rseg
X3266 n_67260_42840 n_67260_45640 Rseg
X3267 n_67260_45640 n_67260_48440 Rseg
X3268 n_67260_48440 n_67260_51240 Rseg
X3269 n_67260_51240 n_67260_54040 Rseg
X3270 n_67260_54040 n_67260_56840 Rseg
X3271 n_67260_56840 n_67260_59640 Rseg
X3272 n_67260_59640 n_67260_62440 Rseg
X3273 n_67260_62440 n_67260_65240 Rseg
X3274 n_67260_65240 n_67260_68040 Rseg
X3275 n_67260_68040 n_67260_70840 Rseg
X3276 n_67260_70840 n_67260_73640 Rseg
X3277 n_67260_73640 n_67260_76440 Rseg
X3278 n_67260_76440 n_67260_79240 Rseg
X3279 n_67260_79240 n_67260_82040 Rseg
X3280 n_67260_82040 n_67260_84840 Rseg
X3281 n_67260_84840 n_67260_87640 Rseg
X3282 n_68020_40040 n_68020_42840 Rseg
X3283 n_68020_42840 n_68020_45640 Rseg
X3284 n_68020_45640 n_68020_48440 Rseg
X3285 n_68020_48440 n_68020_51240 Rseg
X3286 n_68020_51240 n_68020_54040 Rseg
X3287 n_68020_54040 n_68020_56840 Rseg
X3288 n_68020_56840 n_68020_59640 Rseg
X3289 n_68020_59640 n_68020_62440 Rseg
X3290 n_68020_62440 n_68020_65240 Rseg
X3291 n_68020_65240 n_68020_68040 Rseg
X3292 n_68020_68040 n_68020_70840 Rseg
X3293 n_68020_70840 n_68020_73640 Rseg
X3294 n_68020_73640 n_68020_76440 Rseg
X3295 n_68020_76440 n_68020_79240 Rseg
X3296 n_68020_79240 n_68020_82040 Rseg
X3297 n_68020_82040 n_68020_84840 Rseg
X3298 n_68020_84840 n_68020_87640 Rseg
X3299 n_68400_40040 n_68400_42840 Rseg
X3300 n_68400_42840 n_68400_45640 Rseg
X3301 n_68400_45640 n_68400_48440 Rseg
X3302 n_68400_48440 n_68400_51240 Rseg
X3303 n_68400_51240 n_68400_54040 Rseg
X3304 n_68400_54040 n_68400_56840 Rseg
X3305 n_68400_56840 n_68400_59640 Rseg
X3306 n_68400_59640 n_68400_62440 Rseg
X3307 n_68400_62440 n_68400_65240 Rseg
X3308 n_68400_65240 n_68400_68040 Rseg
X3309 n_68400_68040 n_68400_70840 Rseg
X3310 n_68400_70840 n_68400_73640 Rseg
X3311 n_68400_73640 n_68400_76440 Rseg
X3312 n_68400_76440 n_68400_79240 Rseg
X3313 n_68400_79240 n_68400_82040 Rseg
X3314 n_68400_82040 n_68400_84840 Rseg
X3315 n_68400_84840 n_68400_87640 Rseg
X3316 n_68780_40040 n_68780_42840 Rseg
X3317 n_68780_42840 n_68780_45640 Rseg
X3318 n_68780_45640 n_68780_48440 Rseg
X3319 n_68780_48440 n_68780_51240 Rseg
X3320 n_68780_51240 n_68780_54040 Rseg
X3321 n_68780_54040 n_68780_56840 Rseg
X3322 n_68780_56840 n_68780_59640 Rseg
X3323 n_68780_59640 n_68780_62440 Rseg
X3324 n_68780_62440 n_68780_65240 Rseg
X3325 n_68780_65240 n_68780_68040 Rseg
X3326 n_68780_68040 n_68780_70840 Rseg
X3327 n_68780_70840 n_68780_73640 Rseg
X3328 n_68780_73640 n_68780_76440 Rseg
X3329 n_68780_76440 n_68780_79240 Rseg
X3330 n_68780_79240 n_68780_82040 Rseg
X3331 n_68780_82040 n_68780_84840 Rseg
X3332 n_68780_84840 n_68780_87640 Rseg
X3333 n_69160_40040 n_69160_42840 Rseg
X3334 n_69160_42840 n_69160_45640 Rseg
X3335 n_69160_45640 n_69160_48440 Rseg
X3336 n_69160_48440 n_69160_51240 Rseg
X3337 n_69160_51240 n_69160_54040 Rseg
X3338 n_69160_54040 n_69160_56840 Rseg
X3339 n_69160_56840 n_69160_59640 Rseg
X3340 n_69160_59640 n_69160_62440 Rseg
X3341 n_69160_62440 n_69160_65240 Rseg
X3342 n_69160_65240 n_69160_68040 Rseg
X3343 n_69160_68040 n_69160_70840 Rseg
X3344 n_69160_70840 n_69160_73640 Rseg
X3345 n_69160_73640 n_69160_76440 Rseg
X3346 n_69160_76440 n_69160_79240 Rseg
X3347 n_69160_79240 n_69160_82040 Rseg
X3348 n_69160_82040 n_69160_84840 Rseg
X3349 n_69160_84840 n_69160_87640 Rseg
X3350 n_69920_40040 n_69920_42840 Rseg
X3351 n_69920_42840 n_69920_45640 Rseg
X3352 n_69920_45640 n_69920_48440 Rseg
X3353 n_69920_48440 n_69920_51240 Rseg
X3354 n_69920_51240 n_69920_54040 Rseg
X3355 n_69920_54040 n_69920_56840 Rseg
X3356 n_69920_56840 n_69920_59640 Rseg
X3357 n_69920_59640 n_69920_62440 Rseg
X3358 n_69920_62440 n_69920_65240 Rseg
X3359 n_69920_65240 n_69920_68040 Rseg
X3360 n_69920_68040 n_69920_70840 Rseg
X3361 n_69920_70840 n_69920_73640 Rseg
X3362 n_69920_73640 n_69920_76440 Rseg
X3363 n_69920_76440 n_69920_79240 Rseg
X3364 n_69920_79240 n_69920_82040 Rseg
X3365 n_69920_82040 n_69920_84840 Rseg
X3366 n_69920_84840 n_69920_87640 Rseg
X3367 n_70300_40040 n_70300_42840 Rseg
X3368 n_70300_42840 n_70300_45640 Rseg
X3369 n_70300_45640 n_70300_48440 Rseg
X3370 n_70300_48440 n_70300_51240 Rseg
X3371 n_70300_51240 n_70300_54040 Rseg
X3372 n_70300_54040 n_70300_56840 Rseg
X3373 n_70300_56840 n_70300_59640 Rseg
X3374 n_70300_59640 n_70300_62440 Rseg
X3375 n_70300_62440 n_70300_65240 Rseg
X3376 n_70300_65240 n_70300_68040 Rseg
X3377 n_70300_68040 n_70300_70840 Rseg
X3378 n_70300_70840 n_70300_73640 Rseg
X3379 n_70300_73640 n_70300_76440 Rseg
X3380 n_70300_76440 n_70300_79240 Rseg
X3381 n_70300_79240 n_70300_82040 Rseg
X3382 n_70300_82040 n_70300_84840 Rseg
X3383 n_70300_84840 n_70300_87640 Rseg
X3384 n_71060_40040 n_71060_42840 Rseg
X3385 n_71060_42840 n_71060_45640 Rseg
X3386 n_71060_45640 n_71060_48440 Rseg
X3387 n_71060_48440 n_71060_51240 Rseg
X3388 n_71060_51240 n_71060_54040 Rseg
X3389 n_71060_54040 n_71060_56840 Rseg
X3390 n_71060_56840 n_71060_59640 Rseg
X3391 n_71060_59640 n_71060_62440 Rseg
X3392 n_71060_62440 n_71060_65240 Rseg
X3393 n_71060_65240 n_71060_68040 Rseg
X3394 n_71060_68040 n_71060_70840 Rseg
X3395 n_71060_70840 n_71060_73640 Rseg
X3396 n_71060_73640 n_71060_76440 Rseg
X3397 n_71060_76440 n_71060_79240 Rseg
X3398 n_71060_79240 n_71060_82040 Rseg
X3399 n_71060_82040 n_71060_84840 Rseg
X3400 n_71060_84840 n_71060_87640 Rseg
X3401 n_71820_40040 n_71820_42840 Rseg
X3402 n_71820_42840 n_71820_45640 Rseg
X3403 n_71820_45640 n_71820_48440 Rseg
X3404 n_71820_48440 n_71820_51240 Rseg
X3405 n_71820_51240 n_71820_54040 Rseg
X3406 n_71820_54040 n_71820_56840 Rseg
X3407 n_71820_56840 n_71820_59640 Rseg
X3408 n_71820_59640 n_71820_62440 Rseg
X3409 n_71820_62440 n_71820_65240 Rseg
X3410 n_71820_65240 n_71820_68040 Rseg
X3411 n_71820_68040 n_71820_70840 Rseg
X3412 n_71820_70840 n_71820_73640 Rseg
X3413 n_71820_73640 n_71820_76440 Rseg
X3414 n_71820_76440 n_71820_79240 Rseg
X3415 n_71820_79240 n_71820_82040 Rseg
X3416 n_71820_82040 n_71820_84840 Rseg
X3417 n_71820_84840 n_71820_87640 Rseg
X3418 n_72200_40040 n_72200_42840 Rseg
X3419 n_72200_42840 n_72200_45640 Rseg
X3420 n_72200_45640 n_72200_48440 Rseg
X3421 n_72200_48440 n_72200_51240 Rseg
X3422 n_72200_51240 n_72200_54040 Rseg
X3423 n_72200_54040 n_72200_56840 Rseg
X3424 n_72200_56840 n_72200_59640 Rseg
X3425 n_72200_59640 n_72200_62440 Rseg
X3426 n_72200_62440 n_72200_65240 Rseg
X3427 n_72200_65240 n_72200_68040 Rseg
X3428 n_72200_68040 n_72200_70840 Rseg
X3429 n_72200_70840 n_72200_73640 Rseg
X3430 n_72200_73640 n_72200_76440 Rseg
X3431 n_72200_76440 n_72200_79240 Rseg
X3432 n_72200_79240 n_72200_82040 Rseg
X3433 n_72200_82040 n_72200_84840 Rseg
X3434 n_72200_84840 n_72200_87640 Rseg
X3435 n_72960_40040 n_72960_42840 Rseg
X3436 n_72960_42840 n_72960_45640 Rseg
X3437 n_72960_45640 n_72960_48440 Rseg
X3438 n_72960_48440 n_72960_51240 Rseg
X3439 n_72960_51240 n_72960_54040 Rseg
X3440 n_72960_54040 n_72960_56840 Rseg
X3441 n_72960_56840 n_72960_59640 Rseg
X3442 n_72960_59640 n_72960_62440 Rseg
X3443 n_72960_62440 n_72960_65240 Rseg
X3444 n_72960_65240 n_72960_68040 Rseg
X3445 n_72960_68040 n_72960_70840 Rseg
X3446 n_72960_70840 n_72960_73640 Rseg
X3447 n_72960_73640 n_72960_76440 Rseg
X3448 n_72960_76440 n_72960_79240 Rseg
X3449 n_72960_79240 n_72960_82040 Rseg
X3450 n_72960_82040 n_72960_84840 Rseg
X3451 n_72960_84840 n_72960_87640 Rseg
X3452 n_73340_40040 n_73340_42840 Rseg
X3453 n_73340_42840 n_73340_45640 Rseg
X3454 n_73340_45640 n_73340_48440 Rseg
X3455 n_73340_48440 n_73340_51240 Rseg
X3456 n_73340_51240 n_73340_54040 Rseg
X3457 n_73340_54040 n_73340_56840 Rseg
X3458 n_73340_56840 n_73340_59640 Rseg
X3459 n_73340_59640 n_73340_62440 Rseg
X3460 n_73340_62440 n_73340_65240 Rseg
X3461 n_73340_65240 n_73340_68040 Rseg
X3462 n_73340_68040 n_73340_70840 Rseg
X3463 n_73340_70840 n_73340_73640 Rseg
X3464 n_73340_73640 n_73340_76440 Rseg
X3465 n_73340_76440 n_73340_79240 Rseg
X3466 n_73340_79240 n_73340_82040 Rseg
X3467 n_73340_82040 n_73340_84840 Rseg
X3468 n_73340_84840 n_73340_87640 Rseg
X3469 n_73720_40040 n_73720_42840 Rseg
X3470 n_73720_42840 n_73720_45640 Rseg
X3471 n_73720_45640 n_73720_48440 Rseg
X3472 n_73720_48440 n_73720_51240 Rseg
X3473 n_73720_51240 n_73720_54040 Rseg
X3474 n_73720_54040 n_73720_56840 Rseg
X3475 n_73720_56840 n_73720_59640 Rseg
X3476 n_73720_59640 n_73720_62440 Rseg
X3477 n_73720_62440 n_73720_65240 Rseg
X3478 n_73720_65240 n_73720_68040 Rseg
X3479 n_73720_68040 n_73720_70840 Rseg
X3480 n_73720_70840 n_73720_73640 Rseg
X3481 n_73720_73640 n_73720_76440 Rseg
X3482 n_73720_76440 n_73720_79240 Rseg
X3483 n_73720_79240 n_73720_82040 Rseg
X3484 n_73720_82040 n_73720_84840 Rseg
X3485 n_73720_84840 n_73720_87640 Rseg
X3486 n_74100_40040 n_74100_42840 Rseg
X3487 n_74100_42840 n_74100_45640 Rseg
X3488 n_74100_45640 n_74100_48440 Rseg
X3489 n_74100_48440 n_74100_51240 Rseg
X3490 n_74100_51240 n_74100_54040 Rseg
X3491 n_74100_54040 n_74100_56840 Rseg
X3492 n_74100_56840 n_74100_59640 Rseg
X3493 n_74100_59640 n_74100_62440 Rseg
X3494 n_74100_62440 n_74100_65240 Rseg
X3495 n_74100_65240 n_74100_68040 Rseg
X3496 n_74100_68040 n_74100_70840 Rseg
X3497 n_74100_70840 n_74100_73640 Rseg
X3498 n_74100_73640 n_74100_76440 Rseg
X3499 n_74100_76440 n_74100_79240 Rseg
X3500 n_74100_79240 n_74100_82040 Rseg
X3501 n_74100_82040 n_74100_84840 Rseg
X3502 n_74100_84840 n_74100_87640 Rseg
X3503 n_74860_40040 n_74860_42840 Rseg
X3504 n_74860_42840 n_74860_45640 Rseg
X3505 n_74860_45640 n_74860_48440 Rseg
X3506 n_74860_48440 n_74860_51240 Rseg
X3507 n_74860_51240 n_74860_54040 Rseg
X3508 n_74860_54040 n_74860_56840 Rseg
X3509 n_74860_56840 n_74860_59640 Rseg
X3510 n_74860_59640 n_74860_62440 Rseg
X3511 n_74860_62440 n_74860_65240 Rseg
X3512 n_74860_65240 n_74860_68040 Rseg
X3513 n_74860_68040 n_74860_70840 Rseg
X3514 n_74860_70840 n_74860_73640 Rseg
X3515 n_74860_73640 n_74860_76440 Rseg
X3516 n_74860_76440 n_74860_79240 Rseg
X3517 n_74860_79240 n_74860_82040 Rseg
X3518 n_74860_82040 n_74860_84840 Rseg
X3519 n_74860_84840 n_74860_87640 Rseg
X3520 n_75240_40040 n_75240_42840 Rseg
X3521 n_75240_42840 n_75240_45640 Rseg
X3522 n_75240_45640 n_75240_48440 Rseg
X3523 n_75240_48440 n_75240_51240 Rseg
X3524 n_75240_51240 n_75240_54040 Rseg
X3525 n_75240_54040 n_75240_56840 Rseg
X3526 n_75240_56840 n_75240_59640 Rseg
X3527 n_75240_59640 n_75240_62440 Rseg
X3528 n_75240_62440 n_75240_65240 Rseg
X3529 n_75240_65240 n_75240_68040 Rseg
X3530 n_75240_68040 n_75240_70840 Rseg
X3531 n_75240_70840 n_75240_73640 Rseg
X3532 n_75240_73640 n_75240_76440 Rseg
X3533 n_75240_76440 n_75240_79240 Rseg
X3534 n_75240_79240 n_75240_82040 Rseg
X3535 n_75240_82040 n_75240_84840 Rseg
X3536 n_75240_84840 n_75240_87640 Rseg
X3537 n_76000_40040 n_76000_42840 Rseg
X3538 n_76000_42840 n_76000_45640 Rseg
X3539 n_76000_45640 n_76000_48440 Rseg
X3540 n_76000_48440 n_76000_51240 Rseg
X3541 n_76000_51240 n_76000_54040 Rseg
X3542 n_76000_54040 n_76000_56840 Rseg
X3543 n_76000_56840 n_76000_59640 Rseg
X3544 n_76000_59640 n_76000_62440 Rseg
X3545 n_76000_62440 n_76000_65240 Rseg
X3546 n_76000_65240 n_76000_68040 Rseg
X3547 n_76000_68040 n_76000_70840 Rseg
X3548 n_76000_70840 n_76000_73640 Rseg
X3549 n_76000_73640 n_76000_76440 Rseg
X3550 n_76000_76440 n_76000_79240 Rseg
X3551 n_76000_79240 n_76000_82040 Rseg
X3552 n_76000_82040 n_76000_84840 Rseg
X3553 n_76000_84840 n_76000_87640 Rseg
X3554 n_76380_40040 n_76380_42840 Rseg
X3555 n_76380_42840 n_76380_45640 Rseg
X3556 n_76380_45640 n_76380_48440 Rseg
X3557 n_76380_48440 n_76380_51240 Rseg
X3558 n_76380_51240 n_76380_54040 Rseg
X3559 n_76380_54040 n_76380_56840 Rseg
X3560 n_76380_56840 n_76380_59640 Rseg
X3561 n_76380_59640 n_76380_62440 Rseg
X3562 n_76380_62440 n_76380_65240 Rseg
X3563 n_76380_65240 n_76380_68040 Rseg
X3564 n_76380_68040 n_76380_70840 Rseg
X3565 n_76380_70840 n_76380_73640 Rseg
X3566 n_76380_73640 n_76380_76440 Rseg
X3567 n_76380_76440 n_76380_79240 Rseg
X3568 n_76380_79240 n_76380_82040 Rseg
X3569 n_76380_82040 n_76380_84840 Rseg
X3570 n_76380_84840 n_76380_87640 Rseg
X3571 n_76760_40040 n_76760_42840 Rseg
X3572 n_76760_42840 n_76760_45640 Rseg
X3573 n_76760_45640 n_76760_48440 Rseg
X3574 n_76760_48440 n_76760_51240 Rseg
X3575 n_76760_51240 n_76760_54040 Rseg
X3576 n_76760_54040 n_76760_56840 Rseg
X3577 n_76760_56840 n_76760_59640 Rseg
X3578 n_76760_59640 n_76760_62440 Rseg
X3579 n_76760_62440 n_76760_65240 Rseg
X3580 n_76760_65240 n_76760_68040 Rseg
X3581 n_76760_68040 n_76760_70840 Rseg
X3582 n_76760_70840 n_76760_73640 Rseg
X3583 n_76760_73640 n_76760_76440 Rseg
X3584 n_76760_76440 n_76760_79240 Rseg
X3585 n_76760_79240 n_76760_82040 Rseg
X3586 n_76760_82040 n_76760_84840 Rseg
X3587 n_76760_84840 n_76760_87640 Rseg
X3588 n_77140_40040 n_77140_42840 Rseg
X3589 n_77140_42840 n_77140_45640 Rseg
X3590 n_77140_45640 n_77140_48440 Rseg
X3591 n_77140_48440 n_77140_51240 Rseg
X3592 n_77140_51240 n_77140_54040 Rseg
X3593 n_77140_54040 n_77140_56840 Rseg
X3594 n_77140_56840 n_77140_59640 Rseg
X3595 n_77140_59640 n_77140_62440 Rseg
X3596 n_77140_62440 n_77140_65240 Rseg
X3597 n_77140_65240 n_77140_68040 Rseg
X3598 n_77140_68040 n_77140_70840 Rseg
X3599 n_77140_70840 n_77140_73640 Rseg
X3600 n_77140_73640 n_77140_76440 Rseg
X3601 n_77140_76440 n_77140_79240 Rseg
X3602 n_77140_79240 n_77140_82040 Rseg
X3603 n_77140_82040 n_77140_84840 Rseg
X3604 n_77140_84840 n_77140_87640 Rseg
X3605 n_77520_40040 n_77520_42840 Rseg
X3606 n_77520_42840 n_77520_45640 Rseg
X3607 n_77520_45640 n_77520_48440 Rseg
X3608 n_77520_48440 n_77520_51240 Rseg
X3609 n_77520_51240 n_77520_54040 Rseg
X3610 n_77520_54040 n_77520_56840 Rseg
X3611 n_77520_56840 n_77520_59640 Rseg
X3612 n_77520_59640 n_77520_62440 Rseg
X3613 n_77520_62440 n_77520_65240 Rseg
X3614 n_77520_65240 n_77520_68040 Rseg
X3615 n_77520_68040 n_77520_70840 Rseg
X3616 n_77520_70840 n_77520_73640 Rseg
X3617 n_77520_73640 n_77520_76440 Rseg
X3618 n_77520_76440 n_77520_79240 Rseg
X3619 n_77520_79240 n_77520_82040 Rseg
X3620 n_77520_82040 n_77520_84840 Rseg
X3621 n_77520_84840 n_77520_87640 Rseg
X3622 n_77900_40040 n_77900_42840 Rseg
X3623 n_77900_42840 n_77900_45640 Rseg
X3624 n_77900_45640 n_77900_48440 Rseg
X3625 n_77900_48440 n_77900_51240 Rseg
X3626 n_77900_51240 n_77900_54040 Rseg
X3627 n_77900_54040 n_77900_56840 Rseg
X3628 n_77900_56840 n_77900_59640 Rseg
X3629 n_77900_59640 n_77900_62440 Rseg
X3630 n_77900_62440 n_77900_65240 Rseg
X3631 n_77900_65240 n_77900_68040 Rseg
X3632 n_77900_68040 n_77900_70840 Rseg
X3633 n_77900_70840 n_77900_73640 Rseg
X3634 n_77900_73640 n_77900_76440 Rseg
X3635 n_77900_76440 n_77900_79240 Rseg
X3636 n_77900_79240 n_77900_82040 Rseg
X3637 n_77900_82040 n_77900_84840 Rseg
X3638 n_77900_84840 n_77900_87640 Rseg
X3639 n_78280_40040 n_78280_42840 Rseg
X3640 n_78280_42840 n_78280_45640 Rseg
X3641 n_78280_45640 n_78280_48440 Rseg
X3642 n_78280_48440 n_78280_51240 Rseg
X3643 n_78280_51240 n_78280_54040 Rseg
X3644 n_78280_54040 n_78280_56840 Rseg
X3645 n_78280_56840 n_78280_59640 Rseg
X3646 n_78280_59640 n_78280_62440 Rseg
X3647 n_78280_62440 n_78280_65240 Rseg
X3648 n_78280_65240 n_78280_68040 Rseg
X3649 n_78280_68040 n_78280_70840 Rseg
X3650 n_78280_70840 n_78280_73640 Rseg
X3651 n_78280_73640 n_78280_76440 Rseg
X3652 n_78280_76440 n_78280_79240 Rseg
X3653 n_78280_79240 n_78280_82040 Rseg
X3654 n_78280_82040 n_78280_84840 Rseg
X3655 n_78280_84840 n_78280_87640 Rseg
X3656 n_78660_40040 n_78660_42840 Rseg
X3657 n_78660_42840 n_78660_45640 Rseg
X3658 n_78660_45640 n_78660_48440 Rseg
X3659 n_78660_48440 n_78660_51240 Rseg
X3660 n_78660_51240 n_78660_54040 Rseg
X3661 n_78660_54040 n_78660_56840 Rseg
X3662 n_78660_56840 n_78660_59640 Rseg
X3663 n_78660_59640 n_78660_62440 Rseg
X3664 n_78660_62440 n_78660_65240 Rseg
X3665 n_78660_65240 n_78660_68040 Rseg
X3666 n_78660_68040 n_78660_70840 Rseg
X3667 n_78660_70840 n_78660_73640 Rseg
X3668 n_78660_73640 n_78660_76440 Rseg
X3669 n_78660_76440 n_78660_79240 Rseg
X3670 n_78660_79240 n_78660_82040 Rseg
X3671 n_78660_82040 n_78660_84840 Rseg
X3672 n_78660_84840 n_78660_87640 Rseg
X3673 n_79040_40040 n_79040_42840 Rseg
X3674 n_79040_42840 n_79040_45640 Rseg
X3675 n_79040_45640 n_79040_48440 Rseg
X3676 n_79040_48440 n_79040_51240 Rseg
X3677 n_79040_51240 n_79040_54040 Rseg
X3678 n_79040_54040 n_79040_56840 Rseg
X3679 n_79040_56840 n_79040_59640 Rseg
X3680 n_79040_59640 n_79040_62440 Rseg
X3681 n_79040_62440 n_79040_65240 Rseg
X3682 n_79040_65240 n_79040_68040 Rseg
X3683 n_79040_68040 n_79040_70840 Rseg
X3684 n_79040_70840 n_79040_73640 Rseg
X3685 n_79040_73640 n_79040_76440 Rseg
X3686 n_79040_76440 n_79040_79240 Rseg
X3687 n_79040_79240 n_79040_82040 Rseg
X3688 n_79040_82040 n_79040_84840 Rseg
X3689 n_79040_84840 n_79040_87640 Rseg
X3690 n_80180_40040 n_80180_42840 Rseg
X3691 n_80180_42840 n_80180_45640 Rseg
X3692 n_80180_45640 n_80180_48440 Rseg
X3693 n_80180_48440 n_80180_51240 Rseg
X3694 n_80180_51240 n_80180_54040 Rseg
X3695 n_80180_54040 n_80180_56840 Rseg
X3696 n_80180_56840 n_80180_59640 Rseg
X3697 n_80180_59640 n_80180_62440 Rseg
X3698 n_80180_62440 n_80180_65240 Rseg
X3699 n_80180_65240 n_80180_68040 Rseg
X3700 n_80180_68040 n_80180_70840 Rseg
X3701 n_80180_70840 n_80180_73640 Rseg
X3702 n_80180_73640 n_80180_76440 Rseg
X3703 n_80180_76440 n_80180_79240 Rseg
X3704 n_80180_79240 n_80180_82040 Rseg
X3705 n_80180_82040 n_80180_84840 Rseg
X3706 n_80180_84840 n_80180_87640 Rseg
X3707 n_80560_40040 n_80560_42840 Rseg
X3708 n_80560_42840 n_80560_45640 Rseg
X3709 n_80560_45640 n_80560_48440 Rseg
X3710 n_80560_48440 n_80560_51240 Rseg
X3711 n_80560_51240 n_80560_54040 Rseg
X3712 n_80560_54040 n_80560_56840 Rseg
X3713 n_80560_56840 n_80560_59640 Rseg
X3714 n_80560_59640 n_80560_62440 Rseg
X3715 n_80560_62440 n_80560_65240 Rseg
X3716 n_80560_65240 n_80560_68040 Rseg
X3717 n_80560_68040 n_80560_70840 Rseg
X3718 n_80560_70840 n_80560_73640 Rseg
X3719 n_80560_73640 n_80560_76440 Rseg
X3720 n_80560_76440 n_80560_79240 Rseg
X3721 n_80560_79240 n_80560_82040 Rseg
X3722 n_80560_82040 n_80560_84840 Rseg
X3723 n_80560_84840 n_80560_87640 Rseg
X3724 n_80940_40040 n_80940_42840 Rseg
X3725 n_80940_42840 n_80940_45640 Rseg
X3726 n_80940_45640 n_80940_48440 Rseg
X3727 n_80940_48440 n_80940_51240 Rseg
X3728 n_80940_51240 n_80940_54040 Rseg
X3729 n_80940_54040 n_80940_56840 Rseg
X3730 n_80940_56840 n_80940_59640 Rseg
X3731 n_80940_59640 n_80940_62440 Rseg
X3732 n_80940_62440 n_80940_65240 Rseg
X3733 n_80940_65240 n_80940_68040 Rseg
X3734 n_80940_68040 n_80940_70840 Rseg
X3735 n_80940_70840 n_80940_73640 Rseg
X3736 n_80940_73640 n_80940_76440 Rseg
X3737 n_80940_76440 n_80940_79240 Rseg
X3738 n_80940_79240 n_80940_82040 Rseg
X3739 n_80940_82040 n_80940_84840 Rseg
X3740 n_80940_84840 n_80940_87640 Rseg
X3741 n_81700_40040 n_81700_42840 Rseg
X3742 n_81700_42840 n_81700_45640 Rseg
X3743 n_81700_45640 n_81700_48440 Rseg
X3744 n_81700_48440 n_81700_51240 Rseg
X3745 n_81700_51240 n_81700_54040 Rseg
X3746 n_81700_54040 n_81700_56840 Rseg
X3747 n_81700_56840 n_81700_59640 Rseg
X3748 n_81700_59640 n_81700_62440 Rseg
X3749 n_81700_62440 n_81700_65240 Rseg
X3750 n_81700_65240 n_81700_68040 Rseg
X3751 n_81700_68040 n_81700_70840 Rseg
X3752 n_81700_70840 n_81700_73640 Rseg
X3753 n_81700_73640 n_81700_76440 Rseg
X3754 n_81700_76440 n_81700_79240 Rseg
X3755 n_81700_79240 n_81700_82040 Rseg
X3756 n_81700_82040 n_81700_84840 Rseg
X3757 n_81700_84840 n_81700_87640 Rseg
X3758 n_82080_40040 n_82080_42840 Rseg
X3759 n_82080_42840 n_82080_45640 Rseg
X3760 n_82080_45640 n_82080_48440 Rseg
X3761 n_82080_48440 n_82080_51240 Rseg
X3762 n_82080_51240 n_82080_54040 Rseg
X3763 n_82080_54040 n_82080_56840 Rseg
X3764 n_82080_56840 n_82080_59640 Rseg
X3765 n_82080_59640 n_82080_62440 Rseg
X3766 n_82080_62440 n_82080_65240 Rseg
X3767 n_82080_65240 n_82080_68040 Rseg
X3768 n_82080_68040 n_82080_70840 Rseg
X3769 n_82080_70840 n_82080_73640 Rseg
X3770 n_82080_73640 n_82080_76440 Rseg
X3771 n_82080_76440 n_82080_79240 Rseg
X3772 n_82080_79240 n_82080_82040 Rseg
X3773 n_82080_82040 n_82080_84840 Rseg
X3774 n_82080_84840 n_82080_87640 Rseg
X3775 n_83220_40040 n_83220_42840 Rseg
X3776 n_83220_42840 n_83220_45640 Rseg
X3777 n_83220_45640 n_83220_48440 Rseg
X3778 n_83220_48440 n_83220_51240 Rseg
X3779 n_83220_51240 n_83220_54040 Rseg
X3780 n_83220_54040 n_83220_56840 Rseg
X3781 n_83220_56840 n_83220_59640 Rseg
X3782 n_83220_59640 n_83220_62440 Rseg
X3783 n_83220_62440 n_83220_65240 Rseg
X3784 n_83220_65240 n_83220_68040 Rseg
X3785 n_83220_68040 n_83220_70840 Rseg
X3786 n_83220_70840 n_83220_73640 Rseg
X3787 n_83220_73640 n_83220_76440 Rseg
X3788 n_83220_76440 n_83220_79240 Rseg
X3789 n_83220_79240 n_83220_82040 Rseg
X3790 n_83220_82040 n_83220_84840 Rseg
X3791 n_83220_84840 n_83220_87640 Rseg
X3792 n_83600_40040 n_83600_42840 Rseg
X3793 n_83600_42840 n_83600_45640 Rseg
X3794 n_83600_45640 n_83600_48440 Rseg
X3795 n_83600_48440 n_83600_51240 Rseg
X3796 n_83600_51240 n_83600_54040 Rseg
X3797 n_83600_54040 n_83600_56840 Rseg
X3798 n_83600_56840 n_83600_59640 Rseg
X3799 n_83600_59640 n_83600_62440 Rseg
X3800 n_83600_62440 n_83600_65240 Rseg
X3801 n_83600_65240 n_83600_68040 Rseg
X3802 n_83600_68040 n_83600_70840 Rseg
X3803 n_83600_70840 n_83600_73640 Rseg
X3804 n_83600_73640 n_83600_76440 Rseg
X3805 n_83600_76440 n_83600_79240 Rseg
X3806 n_83600_79240 n_83600_82040 Rseg
X3807 n_83600_82040 n_83600_84840 Rseg
X3808 n_83600_84840 n_83600_87640 Rseg
X3809 n_84740_40040 n_84740_42840 Rseg
X3810 n_84740_42840 n_84740_45640 Rseg
X3811 n_84740_45640 n_84740_48440 Rseg
X3812 n_84740_48440 n_84740_51240 Rseg
X3813 n_84740_51240 n_84740_54040 Rseg
X3814 n_84740_54040 n_84740_56840 Rseg
X3815 n_84740_56840 n_84740_59640 Rseg
X3816 n_84740_59640 n_84740_62440 Rseg
X3817 n_84740_62440 n_84740_65240 Rseg
X3818 n_84740_65240 n_84740_68040 Rseg
X3819 n_84740_68040 n_84740_70840 Rseg
X3820 n_84740_70840 n_84740_73640 Rseg
X3821 n_84740_73640 n_84740_76440 Rseg
X3822 n_84740_76440 n_84740_79240 Rseg
X3823 n_84740_79240 n_84740_82040 Rseg
X3824 n_84740_82040 n_84740_84840 Rseg
X3825 n_84740_84840 n_84740_87640 Rseg
X3826 n_85120_40040 n_85120_42840 Rseg
X3827 n_85120_42840 n_85120_45640 Rseg
X3828 n_85120_45640 n_85120_48440 Rseg
X3829 n_85120_48440 n_85120_51240 Rseg
X3830 n_85120_51240 n_85120_54040 Rseg
X3831 n_85120_54040 n_85120_56840 Rseg
X3832 n_85120_56840 n_85120_59640 Rseg
X3833 n_85120_59640 n_85120_62440 Rseg
X3834 n_85120_62440 n_85120_65240 Rseg
X3835 n_85120_65240 n_85120_68040 Rseg
X3836 n_85120_68040 n_85120_70840 Rseg
X3837 n_85120_70840 n_85120_73640 Rseg
X3838 n_85120_73640 n_85120_76440 Rseg
X3839 n_85120_76440 n_85120_79240 Rseg
X3840 n_85120_79240 n_85120_82040 Rseg
X3841 n_85120_82040 n_85120_84840 Rseg
X3842 n_85120_84840 n_85120_87640 Rseg
X3843 n_85500_40040 n_85500_42840 Rseg
X3844 n_85500_42840 n_85500_45640 Rseg
X3845 n_85500_45640 n_85500_48440 Rseg
X3846 n_85500_48440 n_85500_51240 Rseg
X3847 n_85500_51240 n_85500_54040 Rseg
X3848 n_85500_54040 n_85500_56840 Rseg
X3849 n_85500_56840 n_85500_59640 Rseg
X3850 n_85500_59640 n_85500_62440 Rseg
X3851 n_85500_62440 n_85500_65240 Rseg
X3852 n_85500_65240 n_85500_68040 Rseg
X3853 n_85500_68040 n_85500_70840 Rseg
X3854 n_85500_70840 n_85500_73640 Rseg
X3855 n_85500_73640 n_85500_76440 Rseg
X3856 n_85500_76440 n_85500_79240 Rseg
X3857 n_85500_79240 n_85500_82040 Rseg
X3858 n_85500_82040 n_85500_84840 Rseg
X3859 n_85500_84840 n_85500_87640 Rseg
X3860 n_85880_40040 n_85880_42840 Rseg
X3861 n_85880_42840 n_85880_45640 Rseg
X3862 n_85880_45640 n_85880_48440 Rseg
X3863 n_85880_48440 n_85880_51240 Rseg
X3864 n_85880_51240 n_85880_54040 Rseg
X3865 n_85880_54040 n_85880_56840 Rseg
X3866 n_85880_56840 n_85880_59640 Rseg
X3867 n_85880_59640 n_85880_62440 Rseg
X3868 n_85880_62440 n_85880_65240 Rseg
X3869 n_85880_65240 n_85880_68040 Rseg
X3870 n_85880_68040 n_85880_70840 Rseg
X3871 n_85880_70840 n_85880_73640 Rseg
X3872 n_85880_73640 n_85880_76440 Rseg
X3873 n_85880_76440 n_85880_79240 Rseg
X3874 n_85880_79240 n_85880_82040 Rseg
X3875 n_85880_82040 n_85880_84840 Rseg
X3876 n_85880_84840 n_85880_87640 Rseg
X3877 n_86260_40040 n_86260_42840 Rseg
X3878 n_86260_42840 n_86260_45640 Rseg
X3879 n_86260_45640 n_86260_48440 Rseg
X3880 n_86260_48440 n_86260_51240 Rseg
X3881 n_86260_51240 n_86260_54040 Rseg
X3882 n_86260_54040 n_86260_56840 Rseg
X3883 n_86260_56840 n_86260_59640 Rseg
X3884 n_86260_59640 n_86260_62440 Rseg
X3885 n_86260_62440 n_86260_65240 Rseg
X3886 n_86260_65240 n_86260_68040 Rseg
X3887 n_86260_68040 n_86260_70840 Rseg
X3888 n_86260_70840 n_86260_73640 Rseg
X3889 n_86260_73640 n_86260_76440 Rseg
X3890 n_86260_76440 n_86260_79240 Rseg
X3891 n_86260_79240 n_86260_82040 Rseg
X3892 n_86260_82040 n_86260_84840 Rseg
X3893 n_86260_84840 n_86260_87640 Rseg
X3894 n_87020_40040 n_87020_42840 Rseg
X3895 n_87020_42840 n_87020_45640 Rseg
X3896 n_87020_45640 n_87020_48440 Rseg
X3897 n_87020_48440 n_87020_51240 Rseg
X3898 n_87020_51240 n_87020_54040 Rseg
X3899 n_87020_54040 n_87020_56840 Rseg
X3900 n_87020_56840 n_87020_59640 Rseg
X3901 n_87020_59640 n_87020_62440 Rseg
X3902 n_87020_62440 n_87020_65240 Rseg
X3903 n_87020_65240 n_87020_68040 Rseg
X3904 n_87020_68040 n_87020_70840 Rseg
X3905 n_87020_70840 n_87020_73640 Rseg
X3906 n_87020_73640 n_87020_76440 Rseg
X3907 n_87020_76440 n_87020_79240 Rseg
X3908 n_87020_79240 n_87020_82040 Rseg
X3909 n_87020_82040 n_87020_84840 Rseg
X3910 n_87020_84840 n_87020_87640 Rseg
X3911 n_87400_40040 n_87400_42840 Rseg
X3912 n_87400_42840 n_87400_45640 Rseg
X3913 n_87400_45640 n_87400_48440 Rseg
X3914 n_87400_48440 n_87400_51240 Rseg
X3915 n_87400_51240 n_87400_54040 Rseg
X3916 n_87400_54040 n_87400_56840 Rseg
X3917 n_87400_56840 n_87400_59640 Rseg
X3918 n_87400_59640 n_87400_62440 Rseg
X3919 n_87400_62440 n_87400_65240 Rseg
X3920 n_87400_65240 n_87400_68040 Rseg
X3921 n_87400_68040 n_87400_70840 Rseg
X3922 n_87400_70840 n_87400_73640 Rseg
X3923 n_87400_73640 n_87400_76440 Rseg
X3924 n_87400_76440 n_87400_79240 Rseg
X3925 n_87400_79240 n_87400_82040 Rseg
X3926 n_87400_82040 n_87400_84840 Rseg
X3927 n_87400_84840 n_87400_87640 Rseg
X3928 n_87780_40040 n_87780_42840 Rseg
X3929 n_87780_42840 n_87780_45640 Rseg
X3930 n_87780_45640 n_87780_48440 Rseg
X3931 n_87780_48440 n_87780_51240 Rseg
X3932 n_87780_51240 n_87780_54040 Rseg
X3933 n_87780_54040 n_87780_56840 Rseg
X3934 n_87780_56840 n_87780_59640 Rseg
X3935 n_87780_59640 n_87780_62440 Rseg
X3936 n_87780_62440 n_87780_65240 Rseg
X3937 n_87780_65240 n_87780_68040 Rseg
X3938 n_87780_68040 n_87780_70840 Rseg
X3939 n_87780_70840 n_87780_73640 Rseg
X3940 n_87780_73640 n_87780_76440 Rseg
X3941 n_87780_76440 n_87780_79240 Rseg
X3942 n_87780_79240 n_87780_82040 Rseg
X3943 n_87780_82040 n_87780_84840 Rseg
X3944 n_87780_84840 n_87780_87640 Rseg
X3945 n_88160_40040 n_88160_42840 Rseg
X3946 n_88160_42840 n_88160_45640 Rseg
X3947 n_88160_45640 n_88160_48440 Rseg
X3948 n_88160_48440 n_88160_51240 Rseg
X3949 n_88160_51240 n_88160_54040 Rseg
X3950 n_88160_54040 n_88160_56840 Rseg
X3951 n_88160_56840 n_88160_59640 Rseg
X3952 n_88160_59640 n_88160_62440 Rseg
X3953 n_88160_62440 n_88160_65240 Rseg
X3954 n_88160_65240 n_88160_68040 Rseg
X3955 n_88160_68040 n_88160_70840 Rseg
X3956 n_88160_70840 n_88160_73640 Rseg
X3957 n_88160_73640 n_88160_76440 Rseg
X3958 n_88160_76440 n_88160_79240 Rseg
X3959 n_88160_79240 n_88160_82040 Rseg
X3960 n_88160_82040 n_88160_84840 Rseg
X3961 n_88160_84840 n_88160_87640 Rseg
X3962 n_88540_40040 n_88540_42840 Rseg
X3963 n_88540_42840 n_88540_45640 Rseg
X3964 n_88540_45640 n_88540_48440 Rseg
X3965 n_88540_48440 n_88540_51240 Rseg
X3966 n_88540_51240 n_88540_54040 Rseg
X3967 n_88540_54040 n_88540_56840 Rseg
X3968 n_88540_56840 n_88540_59640 Rseg
X3969 n_88540_59640 n_88540_62440 Rseg
X3970 n_88540_62440 n_88540_65240 Rseg
X3971 n_88540_65240 n_88540_68040 Rseg
X3972 n_88540_68040 n_88540_70840 Rseg
X3973 n_88540_70840 n_88540_73640 Rseg
X3974 n_88540_73640 n_88540_76440 Rseg
X3975 n_88540_76440 n_88540_79240 Rseg
X3976 n_88540_79240 n_88540_82040 Rseg
X3977 n_88540_82040 n_88540_84840 Rseg
X3978 n_88540_84840 n_88540_87640 Rseg
X3979 n_88920_40040 n_88920_42840 Rseg
X3980 n_88920_42840 n_88920_45640 Rseg
X3981 n_88920_45640 n_88920_48440 Rseg
X3982 n_88920_48440 n_88920_51240 Rseg
X3983 n_88920_51240 n_88920_54040 Rseg
X3984 n_88920_54040 n_88920_56840 Rseg
X3985 n_88920_56840 n_88920_59640 Rseg
X3986 n_88920_59640 n_88920_62440 Rseg
X3987 n_88920_62440 n_88920_65240 Rseg
X3988 n_88920_65240 n_88920_68040 Rseg
X3989 n_88920_68040 n_88920_70840 Rseg
X3990 n_88920_70840 n_88920_73640 Rseg
X3991 n_88920_73640 n_88920_76440 Rseg
X3992 n_88920_76440 n_88920_79240 Rseg
X3993 n_88920_79240 n_88920_82040 Rseg
X3994 n_88920_82040 n_88920_84840 Rseg
X3995 n_88920_84840 n_88920_87640 Rseg
X3996 n_89300_40040 n_89300_42840 Rseg
X3997 n_89300_42840 n_89300_45640 Rseg
X3998 n_89300_45640 n_89300_48440 Rseg
X3999 n_89300_48440 n_89300_51240 Rseg
X4000 n_89300_51240 n_89300_54040 Rseg
X4001 n_89300_54040 n_89300_56840 Rseg
X4002 n_89300_56840 n_89300_59640 Rseg
X4003 n_89300_59640 n_89300_62440 Rseg
X4004 n_89300_62440 n_89300_65240 Rseg
X4005 n_89300_65240 n_89300_68040 Rseg
X4006 n_89300_68040 n_89300_70840 Rseg
X4007 n_89300_70840 n_89300_73640 Rseg
X4008 n_89300_73640 n_89300_76440 Rseg
X4009 n_89300_76440 n_89300_79240 Rseg
X4010 n_89300_79240 n_89300_82040 Rseg
X4011 n_89300_82040 n_89300_84840 Rseg
X4012 n_89300_84840 n_89300_87640 Rseg
X4013 n_90060_40040 n_90060_42840 Rseg
X4014 n_90060_42840 n_90060_45640 Rseg
X4015 n_90060_45640 n_90060_48440 Rseg
X4016 n_90060_48440 n_90060_51240 Rseg
X4017 n_90060_51240 n_90060_54040 Rseg
X4018 n_90060_54040 n_90060_56840 Rseg
X4019 n_90060_56840 n_90060_59640 Rseg
X4020 n_90060_59640 n_90060_62440 Rseg
X4021 n_90060_62440 n_90060_65240 Rseg
X4022 n_90060_65240 n_90060_68040 Rseg
X4023 n_90060_68040 n_90060_70840 Rseg
X4024 n_90060_70840 n_90060_73640 Rseg
X4025 n_90060_73640 n_90060_76440 Rseg
X4026 n_90060_76440 n_90060_79240 Rseg
X4027 n_90060_79240 n_90060_82040 Rseg
X4028 n_90060_82040 n_90060_84840 Rseg
X4029 n_90060_84840 n_90060_87640 Rseg
X4030 n_90440_40040 n_90440_42840 Rseg
X4031 n_90440_42840 n_90440_45640 Rseg
X4032 n_90440_45640 n_90440_48440 Rseg
X4033 n_90440_48440 n_90440_51240 Rseg
X4034 n_90440_51240 n_90440_54040 Rseg
X4035 n_90440_54040 n_90440_56840 Rseg
X4036 n_90440_56840 n_90440_59640 Rseg
X4037 n_90440_59640 n_90440_62440 Rseg
X4038 n_90440_62440 n_90440_65240 Rseg
X4039 n_90440_65240 n_90440_68040 Rseg
X4040 n_90440_68040 n_90440_70840 Rseg
X4041 n_90440_70840 n_90440_73640 Rseg
X4042 n_90440_73640 n_90440_76440 Rseg
X4043 n_90440_76440 n_90440_79240 Rseg
X4044 n_90440_79240 n_90440_82040 Rseg
X4045 n_90440_82040 n_90440_84840 Rseg
X4046 n_90440_84840 n_90440_87640 Rseg
X4047 n_90820_40040 n_90820_42840 Rseg
X4048 n_90820_42840 n_90820_45640 Rseg
X4049 n_90820_45640 n_90820_48440 Rseg
X4050 n_90820_48440 n_90820_51240 Rseg
X4051 n_90820_51240 n_90820_54040 Rseg
X4052 n_90820_54040 n_90820_56840 Rseg
X4053 n_90820_56840 n_90820_59640 Rseg
X4054 n_90820_59640 n_90820_62440 Rseg
X4055 n_90820_62440 n_90820_65240 Rseg
X4056 n_90820_65240 n_90820_68040 Rseg
X4057 n_90820_68040 n_90820_70840 Rseg
X4058 n_90820_70840 n_90820_73640 Rseg
X4059 n_90820_73640 n_90820_76440 Rseg
X4060 n_90820_76440 n_90820_79240 Rseg
X4061 n_90820_79240 n_90820_82040 Rseg
X4062 n_90820_82040 n_90820_84840 Rseg
X4063 n_90820_84840 n_90820_87640 Rseg
X4064 n_91200_40040 n_91200_42840 Rseg
X4065 n_91200_42840 n_91200_45640 Rseg
X4066 n_91200_45640 n_91200_48440 Rseg
X4067 n_91200_48440 n_91200_51240 Rseg
X4068 n_91200_51240 n_91200_54040 Rseg
X4069 n_91200_54040 n_91200_56840 Rseg
X4070 n_91200_56840 n_91200_59640 Rseg
X4071 n_91200_59640 n_91200_62440 Rseg
X4072 n_91200_62440 n_91200_65240 Rseg
X4073 n_91200_65240 n_91200_68040 Rseg
X4074 n_91200_68040 n_91200_70840 Rseg
X4075 n_91200_70840 n_91200_73640 Rseg
X4076 n_91200_73640 n_91200_76440 Rseg
X4077 n_91200_76440 n_91200_79240 Rseg
X4078 n_91200_79240 n_91200_82040 Rseg
X4079 n_91200_82040 n_91200_84840 Rseg
X4080 n_91200_84840 n_91200_87640 Rseg
X4081 n_91580_40040 n_91580_42840 Rseg
X4082 n_91580_42840 n_91580_45640 Rseg
X4083 n_91580_45640 n_91580_48440 Rseg
X4084 n_91580_48440 n_91580_51240 Rseg
X4085 n_91580_51240 n_91580_54040 Rseg
X4086 n_91580_54040 n_91580_56840 Rseg
X4087 n_91580_56840 n_91580_59640 Rseg
X4088 n_91580_59640 n_91580_62440 Rseg
X4089 n_91580_62440 n_91580_65240 Rseg
X4090 n_91580_65240 n_91580_68040 Rseg
X4091 n_91580_68040 n_91580_70840 Rseg
X4092 n_91580_70840 n_91580_73640 Rseg
X4093 n_91580_73640 n_91580_76440 Rseg
X4094 n_91580_76440 n_91580_79240 Rseg
X4095 n_91580_79240 n_91580_82040 Rseg
X4096 n_91580_82040 n_91580_84840 Rseg
X4097 n_91580_84840 n_91580_87640 Rseg
X4098 n_91960_40040 n_91960_42840 Rseg
X4099 n_91960_42840 n_91960_45640 Rseg
X4100 n_91960_45640 n_91960_48440 Rseg
X4101 n_91960_48440 n_91960_51240 Rseg
X4102 n_91960_51240 n_91960_54040 Rseg
X4103 n_91960_54040 n_91960_56840 Rseg
X4104 n_91960_56840 n_91960_59640 Rseg
X4105 n_91960_59640 n_91960_62440 Rseg
X4106 n_91960_62440 n_91960_65240 Rseg
X4107 n_91960_65240 n_91960_68040 Rseg
X4108 n_91960_68040 n_91960_70840 Rseg
X4109 n_91960_70840 n_91960_73640 Rseg
X4110 n_91960_73640 n_91960_76440 Rseg
X4111 n_91960_76440 n_91960_79240 Rseg
X4112 n_91960_79240 n_91960_82040 Rseg
X4113 n_91960_82040 n_91960_84840 Rseg
X4114 n_91960_84840 n_91960_87640 Rseg
X4115 n_92340_40040 n_92340_42840 Rseg
X4116 n_92340_42840 n_92340_45640 Rseg
X4117 n_92340_45640 n_92340_48440 Rseg
X4118 n_92340_48440 n_92340_51240 Rseg
X4119 n_92340_51240 n_92340_54040 Rseg
X4120 n_92340_54040 n_92340_56840 Rseg
X4121 n_92340_56840 n_92340_59640 Rseg
X4122 n_92340_59640 n_92340_62440 Rseg
X4123 n_92340_62440 n_92340_65240 Rseg
X4124 n_92340_65240 n_92340_68040 Rseg
X4125 n_92340_68040 n_92340_70840 Rseg
X4126 n_92340_70840 n_92340_73640 Rseg
X4127 n_92340_73640 n_92340_76440 Rseg
X4128 n_92340_76440 n_92340_79240 Rseg
X4129 n_92340_79240 n_92340_82040 Rseg
X4130 n_92340_82040 n_92340_84840 Rseg
X4131 n_92340_84840 n_92340_87640 Rseg
X4132 n_92720_40040 n_92720_42840 Rseg
X4133 n_92720_42840 n_92720_45640 Rseg
X4134 n_92720_45640 n_92720_48440 Rseg
X4135 n_92720_48440 n_92720_51240 Rseg
X4136 n_92720_51240 n_92720_54040 Rseg
X4137 n_92720_54040 n_92720_56840 Rseg
X4138 n_92720_56840 n_92720_59640 Rseg
X4139 n_92720_59640 n_92720_62440 Rseg
X4140 n_92720_62440 n_92720_65240 Rseg
X4141 n_92720_65240 n_92720_68040 Rseg
X4142 n_92720_68040 n_92720_70840 Rseg
X4143 n_92720_70840 n_92720_73640 Rseg
X4144 n_92720_73640 n_92720_76440 Rseg
X4145 n_92720_76440 n_92720_79240 Rseg
X4146 n_92720_79240 n_92720_82040 Rseg
X4147 n_92720_82040 n_92720_84840 Rseg
X4148 n_92720_84840 n_92720_87640 Rseg
X4149 n_93100_40040 n_93100_42840 Rseg
X4150 n_93100_42840 n_93100_45640 Rseg
X4151 n_93100_45640 n_93100_48440 Rseg
X4152 n_93100_48440 n_93100_51240 Rseg
X4153 n_93100_51240 n_93100_54040 Rseg
X4154 n_93100_54040 n_93100_56840 Rseg
X4155 n_93100_56840 n_93100_59640 Rseg
X4156 n_93100_59640 n_93100_62440 Rseg
X4157 n_93100_62440 n_93100_65240 Rseg
X4158 n_93100_65240 n_93100_68040 Rseg
X4159 n_93100_68040 n_93100_70840 Rseg
X4160 n_93100_70840 n_93100_73640 Rseg
X4161 n_93100_73640 n_93100_76440 Rseg
X4162 n_93100_76440 n_93100_79240 Rseg
X4163 n_93100_79240 n_93100_82040 Rseg
X4164 n_93100_82040 n_93100_84840 Rseg
X4165 n_93100_84840 n_93100_87640 Rseg
X4166 n_93480_40040 n_93480_42840 Rseg
X4167 n_93480_42840 n_93480_45640 Rseg
X4168 n_93480_45640 n_93480_48440 Rseg
X4169 n_93480_48440 n_93480_51240 Rseg
X4170 n_93480_51240 n_93480_54040 Rseg
X4171 n_93480_54040 n_93480_56840 Rseg
X4172 n_93480_56840 n_93480_59640 Rseg
X4173 n_93480_59640 n_93480_62440 Rseg
X4174 n_93480_62440 n_93480_65240 Rseg
X4175 n_93480_65240 n_93480_68040 Rseg
X4176 n_93480_68040 n_93480_70840 Rseg
X4177 n_93480_70840 n_93480_73640 Rseg
X4178 n_93480_73640 n_93480_76440 Rseg
X4179 n_93480_76440 n_93480_79240 Rseg
X4180 n_93480_79240 n_93480_82040 Rseg
X4181 n_93480_82040 n_93480_84840 Rseg
X4182 n_93480_84840 n_93480_87640 Rseg
* voltage source is placed at (x_min, y_min)
Vin n_40280_40040 0 DC 1.0

I1 n_93480_62440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I2 n_91200_70840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I3 n_93480_79240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I4 n_93480_56840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I5 n_93480_73640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I6 n_93480_76440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I7 n_84740_87640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I8 n_54720_48440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I9 n_40280_54040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I10 n_40660_56840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I11 n_79040_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I12 n_41800_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I13 n_50920_48440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I14 n_63840_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I15 n_70300_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I16 n_91580_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I17 n_87020_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I18 n_88160_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I19 n_52440_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I20 n_40660_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I21 n_42940_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I22 n_56620_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I23 n_67260_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I24 n_90440_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I25 n_93480_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I26 n_80560_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I27 n_46360_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I28 n_40280_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I29 n_40280_48440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I30 n_60040_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I31 n_72200_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I32 n_79040_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I33 n_82080_48440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I34 n_77140_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I35 n_55100_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I36 n_40660_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I37 n_40660_51240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I38 n_60040_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I39 n_43320_59640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I40 n_44460_68040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I41 n_40660_65240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I42 n_41800_68040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I43 n_46740_65240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I44 n_46740_59640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I45 n_57380_48440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I46 n_44840_51240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I47 n_45220_48440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I48 n_54720_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I49 n_74860_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I50 n_80180_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I51 n_76760_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I52 n_71820_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I53 n_56620_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I54 n_41420_48440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I55 n_41420_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I56 n_49400_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I57 n_80180_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I58 n_88920_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I59 n_83600_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I60 n_66880_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I61 n_57760_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I62 n_44840_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I63 n_43700_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I64 n_51680_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I65 n_83600_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I66 n_87020_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I67 n_92720_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I68 n_68400_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I69 n_63460_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I70 n_51680_48440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I71 n_48260_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I72 n_78280_48440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I73 n_41420_54040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I74 n_47880_54040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I75 n_54720_51240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I76 n_81700_87640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I77 n_90440_76440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I78 n_90440_73640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I79 n_88920_56840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I80 n_91580_79240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I81 n_87400_73640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I82 n_91580_62440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I83 n_68780_79240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I84 n_83220_54040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I85 n_91200_54040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I86 n_92340_56840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I87 n_87400_76440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I88 n_92720_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I89 n_87780_87640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I90 n_88920_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I91 n_83600_51240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I92 n_80560_51240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I93 n_85500_51240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I94 n_84740_54040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I95 n_90820_56840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I96 n_77520_54040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I97 n_87400_79240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I98 n_92340_73640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I99 n_88920_76440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I100 n_81700_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I101 n_79040_54040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I102 n_80560_54040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I103 n_82080_54040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I104 n_80560_56840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I105 n_82080_56840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I106 n_78660_56840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I107 n_83600_56840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I108 n_80940_62440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I109 n_76760_56840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I110 n_76380_68040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I111 n_78660_65240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I112 n_77900_68040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I113 n_76000_70840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I114 n_78280_70840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I115 n_75240_73640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I116 n_73720_79240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I117 n_73720_73640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I118 n_67260_84840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I119 n_67260_87640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I120 n_65740_84840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I121 n_62320_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I122 n_65360_87640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I123 n_70300_87640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I124 n_72200_84840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I125 n_82080_51240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I126 n_85500_56840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I127 n_87400_48440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I128 n_85500_59640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I129 n_84740_65240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I130 n_83600_59640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I131 n_82080_68040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I132 n_82080_70840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I133 n_80560_70840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I134 n_80560_73640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I135 n_81700_76440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I136 n_78660_73640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I137 n_78660_76440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I138 n_78660_79240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I139 n_76760_79240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I140 n_80560_79240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I141 n_78660_84840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I142 n_76380_87640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I143 n_74860_84840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I144 n_74860_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I145 n_76760_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I146 n_70300_51240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I147 n_49780_54040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I148 n_52060_51240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I149 n_79040_51240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I150 n_49400_48440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I151 n_53200_48440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I152 n_65360_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I153 n_70300_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I154 n_92720_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I155 n_90440_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I156 n_85500_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I157 n_50540_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I158 n_45220_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I159 n_46740_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I160 n_61560_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I161 n_68020_48440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I162 n_85500_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I163 n_88920_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I164 n_82080_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I165 n_51300_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I166 n_43320_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I167 n_42940_48440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I168 n_53200_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I169 n_73720_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I170 n_76760_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I171 n_82080_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I172 n_73340_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I173 n_53200_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I174 n_44080_48440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I175 n_43320_51240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I176 n_58140_54040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I177 n_58140_56840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I178 n_58520_59640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I179 n_48640_59640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I180 n_52060_54040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I181 n_48260_65240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I182 n_59660_62440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I183 n_50920_68040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I184 n_57380_59640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I185 n_72200_56840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I186 n_49400_65240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I187 n_56620_65240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I188 n_58520_65240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I189 n_60420_65240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I190 n_73720_62440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I191 n_75240_62440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I192 n_63080_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I193 n_75240_59640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I194 n_77520_62440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I195 n_73340_59640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I196 n_46360_76440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I197 n_40660_76440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I198 n_40660_70840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I199 n_66880_73640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I200 n_58140_79240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I201 n_72960_68040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I202 n_68020_62440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I203 n_68780_70840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I204 n_53580_65240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I205 n_53580_68040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I206 n_49400_70840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I207 n_48260_76440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I208 n_45600_84840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I209 n_48640_79240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I210 n_49400_79240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I211 n_60040_76440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I212 n_71820_73640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I213 n_76760_73640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I214 n_56620_79240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I215 n_52060_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I216 n_67260_70840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I217 n_58140_51240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I218 n_49020_68040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I219 n_46360_68040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I220 n_44840_70840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I221 n_43320_70840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I222 n_41800_70840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I223 n_40280_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I224 n_40280_87640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I225 n_57380_76440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I226 n_80560_76440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I227 n_50920_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I228 n_49400_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I229 n_47120_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I230 n_53580_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I231 n_50160_84840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I232 n_65740_73640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I233 n_70300_76440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I234 n_52060_70840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I235 n_52820_79240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I236 n_45220_59640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I237 n_44080_59640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I238 n_42940_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I239 n_42940_84840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I240 n_40280_84840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I241 n_43320_87640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I242 n_61940_84840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I243 n_63080_84840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I244 n_49400_84840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I245 n_52440_87640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I246 n_64220_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I247 n_50920_87640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I248 n_58140_87640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I249 n_59660_84840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I250 n_61940_87640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I251 n_46360_56840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I252 n_46740_51240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I253 n_41800_65240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I254 n_65360_62440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I255 n_66880_62440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I256 n_45220_87640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I257 n_59280_87640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I258 n_51680_84840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I259 n_54340_76440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I260 n_67260_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I261 n_53580_87640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I262 n_64600_84840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I263 n_56240_76440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I264 n_63460_87640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I265 n_67260_65240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I266 n_63460_62440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I267 n_71820_59640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I268 n_71820_70840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I269 n_67260_76440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I270 n_65740_79240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I271 n_64600_79240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I272 n_57380_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I273 n_58520_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I274 n_59660_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I275 n_56240_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I276 n_87400_62440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I277 n_88920_62440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I278 n_87020_59640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I279 n_84740_68040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I280 n_81700_79240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I281 n_85500_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I282 n_68780_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I283 n_71060_82040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I284 n_45220_56840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I285 n_44460_56840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I286 n_60040_59640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I287 n_92340_54040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I288 n_91200_70840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I289 n_87020_87640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I290 n_93100_87640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I291 n_93480_56840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I292 n_93480_76440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I293 n_93100_84840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I294 n_83600_87640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I295 n_65740_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I296 n_61940_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I297 n_40280_54040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I298 n_44080_54040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I299 n_63840_45640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I300 n_79040_42840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I301 n_93480_54040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I302 n_48640_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I303 n_50920_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I304 n_63840_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I305 n_91580_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I306 n_88160_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I307 n_42940_42840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I308 n_56620_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I309 n_67260_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I310 n_93480_45640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I311 n_46360_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I312 n_40280_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I313 n_40280_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I314 n_79040_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I315 n_82080_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I316 n_77140_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I317 n_60040_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I318 n_50160_59640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I319 n_42180_73640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I320 n_44460_68040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I321 n_45600_68040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I322 n_43320_62440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I323 n_47500_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I324 n_44460_62440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I325 n_47500_68040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I326 n_46740_65240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I327 n_52060_73640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I328 n_51300_59640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I329 n_57380_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I330 n_74860_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I331 n_80180_45640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I332 n_76760_42840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I333 n_41420_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I334 n_41420_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I335 n_49400_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I336 n_88920_45640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I337 n_66880_45640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I338 n_57760_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I339 n_44840_45640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I340 n_83600_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I341 n_92720_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I342 n_63460_42840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I343 n_51680_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I344 n_47880_42840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I345 n_92340_51240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I346 n_78280_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I347 n_64980_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I348 n_49020_51240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I349 n_47880_54040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I350 n_60040_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I351 n_63080_51240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I352 n_80180_87640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I353 n_90820_84840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I354 n_90440_76440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I355 n_88920_56840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I356 n_90060_87640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I357 n_85120_84840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I358 n_87400_73640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I359 n_89300_54040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I360 n_73340_51240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I361 n_71820_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I362 n_73340_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I363 n_87780_54040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I364 n_83220_54040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I365 n_91200_54040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I366 n_87400_76440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I367 n_87780_87640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I368 n_88920_82040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I369 n_83600_84840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I370 n_88920_87640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I371 n_83600_51240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I372 n_80560_51240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I373 n_87400_56840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I374 n_88920_76440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I375 n_89300_84840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I376 n_80560_84840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I377 n_77900_51240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I378 n_76380_54040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I379 n_78660_65240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I380 n_80560_65240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I381 n_77900_68040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I382 n_76000_70840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I383 n_75240_73640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I384 n_75240_76440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I385 n_67260_84840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I386 n_71820_79240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I387 n_88920_79240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I388 n_67260_87640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I389 n_65740_84840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I390 n_62320_82040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I391 n_65360_87640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I392 n_70300_84840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I393 n_73720_82040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I394 n_72200_84840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I395 n_87400_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I396 n_82080_59640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I397 n_82080_65240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I398 n_81700_73640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I399 n_81700_76440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I400 n_78660_79240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I401 n_76760_76440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I402 n_72200_76440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I403 n_76760_79240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I404 n_80560_79240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I405 n_78660_84840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I406 n_76760_82040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I407 n_67260_51240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I408 n_61940_51240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I409 n_49780_54040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I410 n_50920_51240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I411 n_61560_54040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I412 n_63080_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I413 n_76380_51240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I414 n_76760_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I415 n_91960_45640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I416 n_83600_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I417 n_85500_45640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I418 n_46360_42840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I419 n_53200_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I420 n_65360_42840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I421 n_89300_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I422 n_81700_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I423 n_43320_45640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I424 n_57380_42840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I425 n_68780_45640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I426 n_83600_45640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I427 n_53580_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I428 n_41800_45640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I429 n_41800_51240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I430 n_74860_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I431 n_80560_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I432 n_75240_42840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I433 n_58140_54040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I434 n_58140_56840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I435 n_58900_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I436 n_58520_59640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I437 n_52060_54040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I438 n_48260_65240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I439 n_44840_73640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I440 n_50920_68040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I441 n_57380_59640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I442 n_40280_59640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I443 n_72200_56840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I444 n_51680_62440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I445 n_56620_65240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I446 n_58520_65240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I447 n_60420_65240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I448 n_73720_62440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I449 n_63460_68040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I450 n_75240_62440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I451 n_76380_59640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I452 n_75240_59640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I453 n_72200_62440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I454 n_41800_62440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I455 n_69160_62440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I456 n_53580_73640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I457 n_49400_73640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I458 n_55860_68040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I459 n_46740_73640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I460 n_46360_76440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I461 n_48260_73640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I462 n_49780_76440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I463 n_50920_79240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I464 n_58520_68040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I465 n_66880_73640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I466 n_58140_79240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I467 n_63460_70840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I468 n_65360_68040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I469 n_68780_68040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I470 n_68020_62440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I471 n_55480_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I472 n_40280_73640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I473 n_68780_70840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I474 n_46740_62440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I475 n_46740_70840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I476 n_48260_76440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I477 n_45600_84840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I478 n_48640_79240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I479 n_49400_79240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I480 n_60040_76440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I481 n_60040_79240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I482 n_63080_79240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I483 n_52060_82040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I484 n_65740_76440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I485 n_67260_70840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I486 n_58140_51240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I487 n_45220_65240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I488 n_70300_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I489 n_49020_68040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I490 n_63080_76440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I491 n_80560_76440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I492 n_50920_82040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I493 n_54720_84840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I494 n_47120_82040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I495 n_53580_82040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I496 n_50160_84840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I497 n_65740_73640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I498 n_47500_56840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I499 n_52060_70840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I500 n_52820_79240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I501 n_45220_59640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I502 n_41420_87640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I503 n_46740_87640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I504 n_43320_87640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I505 n_61940_84840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I506 n_49400_84840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I507 n_52440_87640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I508 n_64220_82040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I509 n_50920_87640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I510 n_58140_87640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I511 n_59660_84840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I512 n_55100_82040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I513 n_46360_56840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I514 n_46740_51240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I515 n_65360_59640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I516 n_65360_56840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I517 n_63080_54040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I518 n_45220_87640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I519 n_59280_87640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I520 n_51680_84840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I521 n_74860_87640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I522 n_67260_82040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I523 n_53580_87640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I524 n_58520_84840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I525 n_56240_76440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I526 n_57000_87640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I527 n_60040_54040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I528 n_66880_59640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I529 n_68400_65240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I530 n_71820_70840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I531 n_67260_76440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I532 n_65740_79240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I533 n_64600_79240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I534 n_57380_82040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I535 n_58520_82040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I536 n_56240_82040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I537 n_87400_62440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I538 n_87020_59640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I539 n_85880_62440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I540 n_83220_65240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I541 n_84740_62440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I542 n_83220_62440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I543 n_83220_68040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I544 n_83600_70840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I545 n_85500_70840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I546 n_84740_73640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I547 n_83600_76440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I548 n_81700_79240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I549 n_85500_76440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I550 n_85500_79240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I551 n_83600_79240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I552 n_85500_82040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I553 n_68780_82040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I554 n_71060_82040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I555 n_61560_56840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I556 n_45220_56840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I557 n_40280_62440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I558 n_44460_56840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I559 n_60040_56840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I560 n_60040_59640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I561 n_92340_54040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I562 n_90820_68040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I563 n_91200_70840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I564 n_87020_87640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I565 n_93100_87640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I566 n_93480_56840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I567 n_90440_62440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I568 n_93480_68040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I569 n_93480_76440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I570 n_56240_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I571 n_65740_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I572 n_61940_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I573 n_40280_54040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I574 n_40660_56840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I575 n_63840_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I576 n_79040_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I577 n_93480_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I578 n_92340_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I579 n_41800_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I580 n_48640_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I581 n_70300_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I582 n_91580_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I583 n_40660_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I584 n_42940_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I585 n_56620_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I586 n_67260_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I587 n_90440_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I588 n_40280_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I589 n_60040_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I590 n_72200_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I591 n_79040_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I592 n_82080_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I593 n_40660_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I594 n_60040_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I595 n_43320_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I596 n_43320_62440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I597 n_40660_65240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I598 n_47500_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I599 n_41800_68040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I600 n_44460_62440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I601 n_46740_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I602 n_57380_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I603 n_45220_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I604 n_80180_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I605 n_76760_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I606 n_71820_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I607 n_56620_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I608 n_41420_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I609 n_83600_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I610 n_66880_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I611 n_57760_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I612 n_44840_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I613 n_43700_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I614 n_92720_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I615 n_68400_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I616 n_47880_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I617 n_48260_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I618 n_85120_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I619 n_90440_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I620 n_78280_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I621 n_64980_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I622 n_41420_54040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I623 n_47880_54040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I624 n_60040_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I625 n_64600_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I626 n_55100_54040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I627 n_90440_76440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I628 n_92340_65240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I629 n_90820_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I630 n_88920_56840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I631 n_90060_87640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I632 n_85120_84840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I633 n_87400_73640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I634 n_88540_68040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I635 n_89300_54040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I636 n_73340_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I637 n_71820_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I638 n_73340_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I639 n_87780_54040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I640 n_88920_70840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I641 n_87400_70840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I642 n_83600_84840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I643 n_88920_87640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I644 n_85500_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I645 n_84740_54040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I646 n_87400_56840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I647 n_77520_54040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I648 n_87400_79240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I649 n_92720_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I650 n_91960_68040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I651 n_90060_79240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I652 n_89300_84840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I653 n_90820_82040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I654 n_80560_84840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I655 n_77900_87640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I656 n_81700_82040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I657 n_79040_87640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I658 n_79040_54040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I659 n_80560_54040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I660 n_77900_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I661 n_82080_54040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I662 n_76380_54040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I663 n_76380_68040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I664 n_77900_68040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I665 n_76000_70840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I666 n_74860_70840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I667 n_73720_70840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I668 n_73720_79240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I669 n_70300_79240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I670 n_67260_84840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I671 n_67260_87640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I672 n_65740_84840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I673 n_65360_87640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I674 n_68780_87640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I675 n_71820_87640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I676 n_70300_87640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I677 n_70300_84840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I678 n_73720_82040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I679 n_72200_84840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I680 n_82080_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I681 n_85500_56840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I682 n_82080_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I683 n_85500_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I684 n_84740_65240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I685 n_82080_65240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I686 n_82080_68040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I687 n_87400_68040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I688 n_82080_70840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I689 n_77140_70840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I690 n_81700_73640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I691 n_80560_70840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I692 n_80560_73640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I693 n_78660_73640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I694 n_79040_70840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I695 n_76380_87640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I696 n_74860_84840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I697 n_76760_82040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I698 n_60800_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I699 n_67260_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I700 n_71820_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I701 n_71820_54040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I702 n_53580_54040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I703 n_56620_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I704 n_59280_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I705 n_49780_54040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I706 n_47880_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I707 n_50920_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I708 n_52060_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I709 n_70300_54040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I710 n_63080_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I711 n_76380_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I712 n_76760_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I713 n_87400_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I714 n_90820_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I715 n_91960_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I716 n_85500_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I717 n_49400_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I718 n_46360_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I719 n_70300_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I720 n_89300_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I721 n_85500_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I722 n_81700_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I723 n_45220_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I724 n_43320_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I725 n_57380_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I726 n_68780_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I727 n_85500_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I728 n_88920_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I729 n_83600_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I730 n_51300_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I731 n_53580_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I732 n_41800_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I733 n_42940_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I734 n_41800_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I735 n_53200_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I736 n_73720_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I737 n_74860_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I738 n_80560_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I739 n_73340_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I740 n_75240_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I741 n_44080_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I742 n_58140_54040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I743 n_56620_56840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I744 n_61940_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I745 n_48640_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I746 n_52060_54040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I747 n_44840_73640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I748 n_40280_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I749 n_72200_56840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I750 n_51680_62440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I751 n_53580_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I752 n_53580_56840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I753 n_49400_65240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I754 n_61560_65240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I755 n_58520_65240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I756 n_59660_68040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I757 n_60420_65240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I758 n_73720_62440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I759 n_66880_68040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I760 n_60800_68040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I761 n_60040_73640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I762 n_63080_65240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I763 n_75240_62440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I764 n_76380_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I765 n_75240_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I766 n_72200_62440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I767 n_61940_68040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I768 n_59660_70840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I769 n_41800_62440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I770 n_53580_73640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I771 n_55100_70840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I772 n_55100_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I773 n_50920_73640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I774 n_46740_73640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I775 n_46360_76440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I776 n_40660_76440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I777 n_48260_73640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I778 n_40660_70840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I779 n_58520_68040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I780 n_58520_73640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I781 n_70300_73640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I782 n_74100_68040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I783 n_75240_65240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I784 n_55480_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I785 n_40280_73640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I786 n_46740_62440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I787 n_53580_65240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I788 n_56240_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I789 n_48260_76440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I790 n_58520_70840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I791 n_60420_70840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I792 n_71820_73640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I793 n_52060_82040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I794 n_65740_76440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I795 n_45220_65240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I796 n_70300_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I797 n_41800_70840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I798 n_40280_82040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I799 n_44080_84840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I800 n_40280_87640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I801 n_50920_82040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I802 n_53580_82040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I803 n_65740_73640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I804 n_47500_56840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I805 n_52820_79240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I806 n_44080_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I807 n_42940_56840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I808 n_41420_87640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I809 n_46740_87640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I810 n_46740_84840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I811 n_49400_84840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I812 n_49400_87640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I813 n_64220_82040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I814 n_55100_82040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I815 n_41800_65240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I816 n_65360_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I817 n_68780_56840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I818 n_45220_87640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I819 n_51680_84840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I820 n_74860_87640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I821 n_67260_82040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I822 n_73340_87640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I823 n_63460_56840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I824 n_68780_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I825 n_67260_56840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I826 n_66880_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I827 n_70300_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I828 n_70300_56840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I829 n_71820_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I830 n_70300_65240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I831 n_71820_65240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I832 n_71820_68040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I833 n_73720_65240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I834 n_70300_68040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I835 n_68780_76440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I836 n_65740_79240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I837 n_53960_79240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I838 n_59660_82040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I839 n_87400_62440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I840 n_87020_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I841 n_83220_65240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I842 n_84740_73640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I843 n_85880_68040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I844 n_85880_73640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I845 n_83600_82040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I846 n_85500_82040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I847 n_69920_82040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I848 n_71060_82040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I849 n_43320_65240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I850 n_40280_62440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I851 n_44460_56840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I852 n_60040_59640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I853 n_93480_62440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I854 n_91200_70840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I855 n_87020_87640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I856 n_93480_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I857 n_93480_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I858 n_83600_87640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I859 n_84740_87640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I860 n_65740_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I861 n_56240_48440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I862 n_65740_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I863 n_61940_48440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I864 n_40280_54040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I865 n_44080_54040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I866 n_40660_56840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I867 n_79040_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I868 n_93480_54040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I869 n_48640_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I870 n_63840_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I871 n_70300_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I872 n_87020_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I873 n_88160_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I874 n_40660_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I875 n_42940_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I876 n_67260_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I877 n_90440_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I878 n_93480_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I879 n_80560_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I880 n_46360_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I881 n_40280_48440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I882 n_79040_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I883 n_82080_48440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I884 n_77140_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I885 n_55100_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I886 n_40660_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I887 n_60040_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I888 n_50160_59640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I889 n_42180_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I890 n_44460_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I891 n_45600_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I892 n_43320_62440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I893 n_40660_65240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I894 n_41800_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I895 n_44460_62440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I896 n_47500_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I897 n_46740_65240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I898 n_52060_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I899 n_51300_59640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I900 n_57380_48440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I901 n_44840_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I902 n_54720_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I903 n_74860_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I904 n_80180_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I905 n_76760_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I906 n_41420_48440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I907 n_49400_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I908 n_80180_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I909 n_88920_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I910 n_83600_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I911 n_66880_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I912 n_44840_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I913 n_43700_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I914 n_83600_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I915 n_87020_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I916 n_68400_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I917 n_63460_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I918 n_47880_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I919 n_92340_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I920 n_78280_48440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I921 n_41420_54040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I922 n_49020_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I923 n_47880_54040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I924 n_60040_48440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I925 n_64600_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I926 n_55100_54040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I927 n_63080_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I928 n_81700_87640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I929 n_80180_87640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I930 n_90440_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I931 n_92340_65240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I932 n_85120_84840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I933 n_87400_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I934 n_91580_62440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I935 n_92340_56840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I936 n_87400_70840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I937 n_83600_84840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I938 n_85500_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I939 n_91960_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I940 n_92340_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I941 n_77900_87640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I942 n_79040_87640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I943 n_80560_56840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I944 n_82080_56840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I945 n_78660_56840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I946 n_76760_65240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I947 n_76760_56840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I948 n_78660_65240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I949 n_80560_65240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I950 n_76000_70840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I951 n_79040_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I952 n_78280_70840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I953 n_74860_70840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I954 n_73720_70840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I955 n_73720_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I956 n_70300_79240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I957 n_67260_84840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I958 n_67260_87640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I959 n_65360_87640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I960 n_68780_87640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I961 n_71820_87640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I962 n_70300_87640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I963 n_70300_84840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I964 n_73720_82040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I965 n_72200_84840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I966 n_82080_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I967 n_87400_48440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I968 n_83600_59640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I969 n_82080_65240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I970 n_82080_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I971 n_85880_65240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I972 n_87400_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I973 n_82080_70840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I974 n_81700_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I975 n_80560_70840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I976 n_80560_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I977 n_78660_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I978 n_79040_70840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I979 n_78660_79240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I980 n_78280_82040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I981 n_80560_79240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I982 n_76760_84840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I983 n_78660_84840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I984 n_76760_82040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I985 n_60800_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I986 n_53580_54040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I987 n_56620_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I988 n_59280_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I989 n_46360_54040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I990 n_47880_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I991 n_41800_56840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I992 n_79040_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I993 n_90820_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I994 n_51680_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I995 n_65360_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I996 n_70300_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I997 n_90440_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I998 n_85500_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I999 n_45220_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1000 n_46740_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1001 n_68020_48440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1002 n_85500_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1003 n_88920_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1004 n_82080_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1005 n_51300_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1006 n_42940_48440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1007 n_76760_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1008 n_82080_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1009 n_73340_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1010 n_53200_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1011 n_43320_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1012 n_58140_54040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1013 n_56620_56840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1014 n_58900_48440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1015 n_57000_54040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1016 n_48260_65240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1017 n_44840_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1018 n_50920_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1019 n_72200_56840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1020 n_53580_59640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1021 n_53580_56840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1022 n_56620_65240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1023 n_61560_65240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1024 n_59660_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1025 n_66880_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1026 n_60800_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1027 n_60040_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1028 n_63080_65240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1029 n_75240_59640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1030 n_72200_62440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1031 n_61940_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1032 n_59660_70840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1033 n_55100_56840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1034 n_69160_62440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1035 n_55100_70840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1036 n_55100_59640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1037 n_50920_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1038 n_46740_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1039 n_46360_76440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1040 n_40660_76440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1041 n_48260_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1042 n_40660_70840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1043 n_58520_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1044 n_58520_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1045 n_70300_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1046 n_63460_70840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1047 n_65360_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1048 n_68780_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1049 n_68020_62440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1050 n_55480_48440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1051 n_53580_65240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1052 n_56240_59640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1053 n_48260_76440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1054 n_58520_70840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1055 n_60420_70840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1056 n_71820_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1057 n_52060_82040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1058 n_65740_76440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1059 n_58140_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1060 n_70300_48440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1061 n_46360_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1062 n_48260_56840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1063 n_41800_70840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1064 n_40280_82040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1065 n_44080_84840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1066 n_40280_87640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1067 n_50920_82040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1068 n_53580_82040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1069 n_65740_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1070 n_47500_56840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1071 n_52820_79240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1072 n_44080_59640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1073 n_42940_56840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1074 n_41420_87640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1075 n_46740_87640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1076 n_46740_84840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1077 n_49400_84840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1078 n_49400_87640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1079 n_64220_82040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1080 n_55100_82040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1081 n_42940_54040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1082 n_43320_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1083 n_44080_65240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1084 n_63080_54040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1085 n_68780_56840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1086 n_45220_87640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1087 n_51680_84840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1088 n_67260_82040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1089 n_73340_87640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1090 n_63460_56840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1091 n_60040_54040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1092 n_68780_59640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1093 n_67260_56840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1094 n_70300_59640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1095 n_70300_56840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1096 n_70300_65240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1097 n_71820_65240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1098 n_71820_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1099 n_73720_65240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1100 n_70300_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1101 n_68780_76440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1102 n_65740_79240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1103 n_53960_79240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1104 n_59660_82040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1105 n_88160_59640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1106 n_83220_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1107 n_84740_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1108 n_83220_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1109 n_84740_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1110 n_85880_68040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1111 n_85880_73640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1112 n_87400_82040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1113 n_83600_82040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1114 n_69920_82040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1115 n_71060_82040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1116 n_43320_65240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I1117 n_93480_79240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1118 n_93100_87640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1119 n_93480_56840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1120 n_93480_68040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1121 n_93480_73640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1122 n_84740_87640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1123 n_65740_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1124 n_54720_48440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1125 n_56240_48440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1126 n_61940_48440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1127 n_63840_45640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1128 n_92340_48440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1129 n_48640_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1130 n_50920_48440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1131 n_70300_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1132 n_42940_42840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1133 n_56620_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1134 n_67260_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1135 n_93480_45640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1136 n_80560_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1137 n_46360_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1138 n_40280_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1139 n_72200_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1140 n_79040_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1141 n_77140_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1142 n_55100_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1143 n_42180_73640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1144 n_45600_68040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1145 n_47500_68040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1146 n_52060_73640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1147 n_54720_42840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1148 n_74860_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1149 n_76760_42840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1150 n_71820_42840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1151 n_41420_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1152 n_49400_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1153 n_80180_42840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1154 n_88920_45640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1155 n_66880_45640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1156 n_57760_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1157 n_44840_45640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1158 n_68400_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1159 n_51680_48440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1160 n_47880_42840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1161 n_85120_48440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1162 n_64980_48440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1163 n_60040_48440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1164 n_55100_54040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1165 n_54720_51240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1166 n_63080_51240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1167 n_81700_87640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1168 n_90440_73640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1169 n_92340_65240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1170 n_88920_56840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1171 n_90060_87640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1172 n_91580_79240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1173 n_83220_54040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1174 n_91200_54040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1175 n_92340_56840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1176 n_90820_65240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1177 n_88920_70840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1178 n_87400_65240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1179 n_92340_76440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1180 n_87780_87640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1181 n_88920_82040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1182 n_83600_84840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1183 n_82080_84840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1184 n_85880_87640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1185 n_83600_51240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1186 n_80560_51240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1187 n_84740_54040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1188 n_87400_56840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1189 n_77520_54040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1190 n_87400_79240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1191 n_89300_59640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1192 n_92720_59640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1193 n_88920_65240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1194 n_92340_73640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1195 n_88920_76440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1196 n_90060_79240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1197 n_89300_84840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1198 n_90820_82040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1199 n_81700_82040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1200 n_79040_54040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1201 n_80560_54040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1202 n_82080_54040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1203 n_80560_56840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1204 n_80180_59640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1205 n_82080_56840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1206 n_78660_56840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1207 n_76380_54040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1208 n_76760_65240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1209 n_78660_65240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1210 n_77900_68040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1211 n_79040_68040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1212 n_78280_70840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1213 n_75240_76440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1214 n_70300_79240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1215 n_67260_84840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1216 n_67260_87640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1217 n_65360_87640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1218 n_70300_84840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1219 n_73720_82040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1220 n_72200_84840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1221 n_85500_56840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1222 n_86260_54040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1223 n_82080_59640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1224 n_84740_65240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1225 n_83600_59640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1226 n_85880_65240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1227 n_87400_68040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1228 n_80560_70840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1229 n_80560_73640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1230 n_76760_76440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1231 n_72200_76440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1232 n_74860_82040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1233 n_67260_51240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1234 n_71820_51240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1235 n_71820_54040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1236 n_70300_51240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1237 n_68020_54040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1238 n_61940_51240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1239 n_46360_54040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1240 n_49780_54040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1241 n_41800_56840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1242 n_52060_51240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1243 n_70300_54040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1244 n_61560_54040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1245 n_66120_51240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1246 n_83600_48440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1247 n_51680_45640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1248 n_53200_48440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1249 n_70300_42840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1250 n_46740_45640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1251 n_61560_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1252 n_68020_48440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1253 n_88920_42840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1254 n_82080_42840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1255 n_51300_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1256 n_43320_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1257 n_73720_45640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1258 n_76760_45640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1259 n_73340_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1260 n_53200_42840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1261 n_58900_48440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1262 n_57000_54040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1263 n_61940_59640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1264 n_52060_54040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1265 n_48260_65240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1266 n_44840_73640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1267 n_50920_68040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1268 n_56620_65240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1269 n_61560_62440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1270 n_61560_65240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1271 n_59660_68040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1272 n_66880_68040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1273 n_60800_68040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1274 n_60040_73640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1275 n_63080_65240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1276 n_61940_68040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1277 n_59660_70840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1278 n_55100_56840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1279 n_69160_62440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1280 n_55100_70840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1281 n_53580_70840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1282 n_55100_73640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1283 n_50920_73640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1284 n_46740_73640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1285 n_46360_76440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1286 n_40660_76440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1287 n_48260_73640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1288 n_40660_70840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1289 n_58520_68040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1290 n_58520_73640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1291 n_56620_73640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1292 n_58140_79240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1293 n_63460_70840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1294 n_65360_68040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1295 n_68780_68040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1296 n_68020_62440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1297 n_48260_76440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1298 n_47500_79240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1299 n_48640_79240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1300 n_58520_70840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1301 n_60040_76440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1302 n_60420_70840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1303 n_63080_73640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1304 n_60040_79240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1305 n_63080_79240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1306 n_52060_82040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1307 n_65740_76440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1308 n_58140_51240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1309 n_70300_48440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1310 n_46360_68040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1311 n_48260_56840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1312 n_40660_79240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1313 n_40280_82040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1314 n_43700_79240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1315 n_40280_87640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1316 n_63080_76440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1317 n_50920_82040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1318 n_53580_82040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1319 n_65740_73640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1320 n_47500_56840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1321 n_52820_79240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1322 n_40280_84840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1323 n_41420_87640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1324 n_46740_87640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1325 n_46740_84840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1326 n_49400_84840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1327 n_52440_87640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1328 n_49400_87640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1329 n_64220_82040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1330 n_58140_87640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1331 n_55100_82040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1332 n_46740_51240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1333 n_44080_65240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1334 n_43320_76440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1335 n_44080_82040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1336 n_63080_54040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1337 n_68780_56840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1338 n_54340_87640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1339 n_67260_82040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1340 n_53580_87640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1341 n_73340_87640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1342 n_57000_87640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1343 n_65360_65240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1344 n_63460_62440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1345 n_63460_59640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1346 n_63460_56840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1347 n_60040_54040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1348 n_67260_56840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1349 n_70300_59640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1350 n_70300_62440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1351 n_70300_65240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1352 n_71820_65240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1353 n_71820_68040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1354 n_70300_70840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1355 n_70300_68040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1356 n_67260_76440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1357 n_65740_79240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1358 n_53960_79240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1359 n_59660_82040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1360 n_56240_82040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1361 n_83220_65240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1362 n_83220_68040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1363 n_84740_68040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1364 n_83220_73640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1365 n_85880_68040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1366 n_83600_82040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1367 n_69920_82040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1368 n_71060_82040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1369 n_72200_82040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1370 n_61560_56840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1371 n_44460_56840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I1372 n_92340_54040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1373 n_93480_62440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1374 n_90820_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1375 n_91200_70840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1376 n_91960_87640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1377 n_93100_87640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1378 n_93480_56840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1379 n_90440_62440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1380 n_93480_76440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1381 n_93100_84840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1382 n_84740_87640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1383 n_65740_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1384 n_65740_45640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1385 n_61940_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1386 n_40660_56840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1387 n_63840_45640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1388 n_79040_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1389 n_93480_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1390 n_92340_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1391 n_91580_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1392 n_40660_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1393 n_56620_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1394 n_90440_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1395 n_80560_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1396 n_46360_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1397 n_40280_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1398 n_60040_45640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1399 n_72200_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1400 n_82080_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1401 n_77140_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1402 n_55100_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1403 n_60040_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1404 n_42180_73640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1405 n_45600_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1406 n_43320_62440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1407 n_40660_65240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1408 n_47500_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1409 n_89300_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1410 n_41800_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1411 n_44460_62440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1412 n_47500_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1413 n_52060_73640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1414 n_57380_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1415 n_54720_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1416 n_74860_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1417 n_80180_45640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1418 n_71820_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1419 n_56620_45640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1420 n_41420_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1421 n_49400_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1422 n_80180_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1423 n_83600_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1424 n_57760_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1425 n_43700_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1426 n_92720_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1427 n_85120_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1428 n_90440_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1429 n_78280_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1430 n_64980_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1431 n_41420_54040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1432 n_60040_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1433 n_64600_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1434 n_63080_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1435 n_81700_87640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1436 n_90820_84840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1437 n_90440_76440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1438 n_90820_59640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1439 n_88920_56840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1440 n_90060_87640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1441 n_87400_84840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1442 n_87400_73640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1443 n_88540_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1444 n_91580_62440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1445 n_89300_54040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1446 n_73340_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1447 n_71820_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1448 n_73340_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1449 n_73720_54040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1450 n_88920_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1451 n_90820_65240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1452 n_87400_65240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1453 n_87400_76440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1454 n_88920_82040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1455 n_85880_87640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1456 n_83600_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1457 n_80560_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1458 n_84740_54040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1459 n_87400_56840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1460 n_77520_54040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1461 n_87400_79240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1462 n_89300_59640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1463 n_88920_65240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1464 n_91960_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1465 n_88920_76440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1466 n_89300_84840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1467 n_81700_82040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1468 n_79040_54040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1469 n_80560_54040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1470 n_82080_54040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1471 n_82080_56840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1472 n_78660_56840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1473 n_76760_65240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1474 n_80940_62440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1475 n_78660_65240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1476 n_77900_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1477 n_76000_70840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1478 n_75240_73640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1479 n_73720_79240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1480 n_73720_73640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1481 n_70300_79240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1482 n_67260_84840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1483 n_71820_79240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1484 n_88920_79240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1485 n_67260_87640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1486 n_65740_84840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1487 n_65360_87640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1488 n_70300_84840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1489 n_73720_82040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1490 n_72200_84840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1491 n_85500_56840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1492 n_86260_54040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1493 n_87400_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1494 n_82080_59640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1495 n_84740_65240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1496 n_83600_59640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1497 n_82080_65240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1498 n_85880_65240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1499 n_87400_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1500 n_81700_73640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1501 n_80560_70840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1502 n_80560_73640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1503 n_78660_73640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1504 n_78660_76440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1505 n_78660_79240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1506 n_78280_82040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1507 n_80560_79240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1508 n_76760_84840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1509 n_78660_84840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1510 n_76380_87640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1511 n_74860_84840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1512 n_74860_82040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1513 n_67260_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1514 n_71820_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1515 n_71820_54040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1516 n_53200_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1517 n_70300_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1518 n_53580_54040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1519 n_68020_54040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1520 n_56620_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1521 n_61940_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1522 n_46360_54040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1523 n_49780_54040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1524 n_52060_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1525 n_75240_54040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1526 n_66120_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1527 n_76380_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1528 n_79040_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1529 n_87400_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1530 n_83600_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1531 n_49400_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1532 n_50160_45640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1533 n_53200_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1534 n_48260_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1535 n_65360_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1536 n_61560_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1537 n_70300_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1538 n_68020_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1539 n_89300_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1540 n_90440_45640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1541 n_87400_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1542 n_44840_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1543 n_61560_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1544 n_78660_45640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1545 n_88920_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1546 n_83600_45640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1547 n_73720_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1548 n_51300_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1549 n_43320_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1550 n_53200_45640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1551 n_71820_45640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1552 n_82080_45640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1553 n_73340_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1554 n_55100_62440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1555 n_44080_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1556 n_46740_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1557 n_43320_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1558 n_45220_54040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1559 n_60040_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1560 n_57000_54040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1561 n_72200_56840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1562 n_61560_62440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1563 n_61560_65240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1564 n_58520_65240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1565 n_59660_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1566 n_60420_65240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1567 n_73720_62440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1568 n_66880_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1569 n_60800_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1570 n_60040_73640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1571 n_63080_65240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1572 n_75240_62440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1573 n_76380_59640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1574 n_75240_59640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1575 n_72200_62440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1576 n_61940_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1577 n_59660_70840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1578 n_69160_62440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1579 n_55100_70840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1580 n_53580_70840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1581 n_55100_73640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1582 n_46360_76440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1583 n_48260_73640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1584 n_58520_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1585 n_58520_73640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1586 n_56620_73640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1587 n_66880_73640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1588 n_63460_70840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1589 n_65360_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1590 n_68780_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1591 n_68020_62440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1592 n_55480_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1593 n_68780_70840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1594 n_46740_70840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1595 n_48260_76440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1596 n_47500_79240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1597 n_58520_70840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1598 n_60420_70840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1599 n_63080_73640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1600 n_67260_70840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1601 n_58140_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1602 n_49020_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1603 n_44080_84840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1604 n_40280_87640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1605 n_47120_82040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1606 n_50160_84840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1607 n_47500_56840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1608 n_40280_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1609 n_45220_59640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1610 n_41420_87640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1611 n_46740_87640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1612 n_46740_84840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1613 n_49400_87640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1614 n_64220_82040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1615 n_50920_87640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1616 n_59660_84840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1617 n_41800_59640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1618 n_43320_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1619 n_43320_76440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1620 n_44080_82040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1621 n_65360_59640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1622 n_45220_87640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1623 n_59280_87640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1624 n_74860_87640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1625 n_54340_87640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1626 n_67260_82040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1627 n_58520_84840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1628 n_73340_87640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1629 n_56240_76440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1630 n_70300_62440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1631 n_70300_56840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1632 n_70300_65240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1633 n_71820_65240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1634 n_71820_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1635 n_70300_70840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1636 n_70300_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1637 n_71820_70840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1638 n_64600_79240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1639 n_57380_82040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1640 n_58520_82040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1641 n_59660_82040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1642 n_56620_84840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1643 n_87400_62440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1644 n_88920_62440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1645 n_88160_59640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1646 n_85880_62440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1647 n_83220_65240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1648 n_84740_62440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1649 n_83220_62440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1650 n_83220_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1651 n_83600_70840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1652 n_85500_70840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1653 n_84740_73640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1654 n_85880_68040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1655 n_83600_76440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1656 n_85500_76440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1657 n_85500_79240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1658 n_87400_82040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1659 n_83600_82040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1660 n_83600_79240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1661 n_85500_82040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1662 n_69920_82040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1663 n_71060_82040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1664 n_72200_82040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1665 n_43320_65240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1666 n_44460_56840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1667 n_60040_59640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I1668 n_92340_54040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1669 n_93480_79240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1670 n_91960_87640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1671 n_93100_87640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1672 n_93480_76440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1673 n_84740_87640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1674 n_54720_48440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1675 n_56240_48440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1676 n_44080_54040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1677 n_40660_56840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1678 n_93480_54040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1679 n_48640_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1680 n_63840_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1681 n_70300_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1682 n_91580_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1683 n_87020_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1684 n_88160_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1685 n_67260_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1686 n_90440_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1687 n_93480_45640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1688 n_80560_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1689 n_46360_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1690 n_40280_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1691 n_60040_45640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1692 n_79040_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1693 n_82080_48440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1694 n_77140_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1695 n_55100_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1696 n_40660_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1697 n_60040_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1698 n_42180_73640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1699 n_44460_68040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1700 n_43320_62440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1701 n_40660_65240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1702 n_47500_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1703 n_89300_48440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1704 n_41800_68040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1705 n_44460_62440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1706 n_46740_65240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1707 n_52060_73640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1708 n_57380_48440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1709 n_44840_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1710 n_54720_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1711 n_74860_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1712 n_80180_45640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1713 n_76760_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1714 n_56620_45640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1715 n_41420_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1716 n_49400_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1717 n_80180_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1718 n_88920_45640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1719 n_83600_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1720 n_66880_45640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1721 n_83600_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1722 n_87020_45640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1723 n_92720_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1724 n_68400_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1725 n_63460_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1726 n_47880_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1727 n_92340_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1728 n_41420_54040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1729 n_49020_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1730 n_55100_54040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1731 n_54720_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1732 n_81700_87640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1733 n_90440_76440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1734 n_90060_87640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1735 n_87400_84840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1736 n_91580_79240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1737 n_89300_54040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1738 n_73340_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1739 n_71820_48440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1740 n_73340_48440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1741 n_73720_54040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1742 n_88920_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1743 n_83220_54040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1744 n_91200_54040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1745 n_87400_70840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1746 n_87400_76440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1747 n_92340_76440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1748 n_87780_87640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1749 n_83600_84840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1750 n_82080_84840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1751 n_88920_87640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1752 n_80560_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1753 n_85500_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1754 n_84740_54040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1755 n_90060_79240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1756 n_79040_87640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1757 n_80180_59640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1758 n_82080_56840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1759 n_78660_56840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1760 n_76380_54040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1761 n_76760_65240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1762 n_80940_62440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1763 n_76760_56840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1764 n_76380_68040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1765 n_75240_73640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1766 n_74860_70840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1767 n_73720_70840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1768 n_75240_76440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1769 n_71820_79240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1770 n_88920_79240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1771 n_82080_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1772 n_85500_56840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1773 n_85500_59640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1774 n_84740_65240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1775 n_83600_59640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1776 n_85880_65240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1777 n_87400_68040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1778 n_82080_70840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1779 n_80560_68040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1780 n_77140_70840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1781 n_80560_70840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1782 n_80560_73640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1783 n_79040_70840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1784 n_78660_76440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1785 n_76760_76440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1786 n_72200_76440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1787 n_76380_87640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1788 n_74860_84840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1789 n_71820_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1790 n_71820_54040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1791 n_53200_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1792 n_53580_54040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1793 n_56620_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1794 n_68780_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1795 n_46360_54040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1796 n_49780_54040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1797 n_50920_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1798 n_52060_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1799 n_75240_54040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1800 n_76380_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1801 n_90820_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1802 n_49400_48440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1803 n_50160_45640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1804 n_51680_45640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1805 n_53200_48440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1806 n_48260_48440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1807 n_61560_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1808 n_68020_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1809 n_89300_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1810 n_87400_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1811 n_85500_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1812 n_45220_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1813 n_44840_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1814 n_68020_48440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1815 n_78660_45640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1816 n_83600_45640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1817 n_73720_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1818 n_51300_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1819 n_43320_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1820 n_53200_45640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1821 n_73720_45640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1822 n_71820_45640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1823 n_76760_45640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1824 n_82080_45640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1825 n_73340_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1826 n_55100_62440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1827 n_44080_48440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1828 n_46740_48440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1829 n_45220_54040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1830 n_60040_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1831 n_57000_54040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1832 n_72200_56840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1833 n_61560_62440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1834 n_75240_59640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1835 n_77520_62440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1836 n_72200_62440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1837 n_69160_62440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1838 n_55100_70840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1839 n_53580_70840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1840 n_55100_73640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1841 n_61560_73640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1842 n_58520_73640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1843 n_70300_73640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1844 n_58140_79240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1845 n_63460_70840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1846 n_74100_68040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1847 n_65360_68040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1848 n_68780_68040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1849 n_75240_65240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1850 n_68020_62440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1851 n_55480_48440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1852 n_53580_65240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1853 n_53580_68040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1854 n_54720_68040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1855 n_48640_79240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1856 n_60040_76440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1857 n_63080_73640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1858 n_71820_73640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1859 n_60040_79240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1860 n_63080_79240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1861 n_58140_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1862 n_49020_68040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1863 n_46360_68040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1864 n_44840_70840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1865 n_44840_76440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1866 n_41800_70840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1867 n_40660_79240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1868 n_43700_79240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1869 n_40280_87640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1870 n_63080_76440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1871 n_47120_82040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1872 n_53580_82040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1873 n_40280_68040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1874 n_52820_79240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1875 n_45220_59640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1876 n_40280_84840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1877 n_41420_87640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1878 n_46740_87640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1879 n_46740_84840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1880 n_49400_84840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1881 n_55100_82040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1882 n_42940_54040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1883 n_41800_59640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1884 n_43320_68040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1885 n_43320_76440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1886 n_44080_82040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1887 n_65360_59640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1888 n_74860_87640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1889 n_73340_87640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1890 n_70300_59640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1891 n_70300_56840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1892 n_71820_59640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1893 n_71820_70840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1894 n_67260_76440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1895 n_68780_76440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1896 n_53960_79240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1897 n_83220_62440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1898 n_83220_68040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1899 n_83600_70840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1900 n_85500_70840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1901 n_85880_68040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1902 n_85880_73640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1903 n_83600_76440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1904 n_85500_76440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1905 n_85500_79240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1906 n_83600_79240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1907 n_69920_82040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1908 n_71060_82040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1909 n_72200_82040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1910 n_43320_65240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1911 n_60040_59640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I1912 n_90820_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1913 n_93480_79240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1914 n_91960_87640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1915 n_93100_87640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1916 n_93480_73640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1917 n_83600_87640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1918 n_84740_87640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1919 n_56240_48440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1920 n_61940_48440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1921 n_40280_54040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1922 n_40660_56840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1923 n_79040_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1924 n_93480_48440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1925 n_93480_54040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1926 n_92340_48440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1927 n_87020_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1928 n_88160_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1929 n_52440_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1930 n_40660_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1931 n_42940_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1932 n_56620_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1933 n_80560_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1934 n_46360_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1935 n_40280_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1936 n_72200_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1937 n_77140_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1938 n_55100_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1939 n_40660_51240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1940 n_43320_59640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1941 n_44460_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1942 n_47500_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1943 n_46740_65240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1944 n_46740_59640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1945 n_44840_51240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1946 n_54720_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1947 n_74860_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1948 n_71820_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1949 n_41420_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1950 n_49400_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1951 n_80180_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1952 n_57760_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1953 n_44840_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1954 n_43700_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1955 n_51680_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1956 n_83600_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1957 n_87020_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1958 n_85120_48440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1959 n_92340_51240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1960 n_90440_48440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1961 n_78280_48440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1962 n_41420_54040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1963 n_47880_54040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1964 n_60040_48440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1965 n_55100_54040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1966 n_81700_87640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1967 n_80180_87640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1968 n_90440_73640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1969 n_90060_87640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1970 n_87400_84840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1971 n_91580_79240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1972 n_88540_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1973 n_73340_51240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1974 n_71820_48440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1975 n_73340_48440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1976 n_88920_70840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1977 n_92720_82040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1978 n_87780_87640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1979 n_88920_87640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1980 n_80560_51240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1981 n_84740_54040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1982 n_77520_54040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1983 n_87400_79240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1984 n_88920_65240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1985 n_91960_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1986 n_89300_73640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1987 n_88920_76440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1988 n_90060_79240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1989 n_80560_84840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1990 n_79040_87640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1991 n_79040_54040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1992 n_77900_51240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1993 n_80560_56840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1994 n_82080_56840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1995 n_83600_56840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1996 n_76380_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1997 n_78660_65240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1998 n_80560_65240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I1999 n_79040_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2000 n_78280_70840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2001 n_75240_76440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2002 n_73720_79240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2003 n_70300_79240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2004 n_67260_84840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2005 n_67260_87640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2006 n_65740_84840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2007 n_62320_82040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2008 n_68780_87640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2009 n_68780_84840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2010 n_70300_87640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2011 n_70300_84840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2012 n_72200_84840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2013 n_85500_56840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2014 n_85500_59640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2015 n_84740_65240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2016 n_82080_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2017 n_85880_65240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2018 n_87400_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2019 n_80560_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2020 n_77140_70840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2021 n_80560_73640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2022 n_81700_76440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2023 n_79040_70840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2024 n_78660_76440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2025 n_76760_76440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2026 n_72200_76440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2027 n_80180_82040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2028 n_76760_84840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2029 n_78660_84840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2030 n_74860_84840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2031 n_76760_82040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2032 n_68020_54040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2033 n_61940_51240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2034 n_49780_54040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2035 n_52060_51240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2036 n_76380_51240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2037 n_76760_48440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2038 n_90820_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2039 n_90820_51240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2040 n_85500_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2041 n_49400_48440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2042 n_50160_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2043 n_51680_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2044 n_46360_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2045 n_53200_48440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2046 n_48260_48440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2047 n_87400_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2048 n_85500_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2049 n_49400_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2050 n_45220_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2051 n_43320_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2052 n_57380_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2053 n_68020_48440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2054 n_68780_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2055 n_73720_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2056 n_51300_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2057 n_43320_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2058 n_53200_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2059 n_58520_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2060 n_73720_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2061 n_76760_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2062 n_74860_48440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2063 n_82080_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2064 n_80560_48440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2065 n_73340_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2066 n_55100_62440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2067 n_44080_48440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2068 n_46740_48440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2069 n_45220_54040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2070 n_58900_48440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2071 n_57000_54040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2072 n_48640_59640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2073 n_52060_54040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2074 n_48260_65240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2075 n_50920_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2076 n_40280_59640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2077 n_49400_65240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2078 n_56620_65240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2079 n_61560_62440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2080 n_58520_65240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2081 n_59660_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2082 n_66880_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2083 n_60800_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2084 n_60040_73640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2085 n_63080_65240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2086 n_61940_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2087 n_59660_70840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2088 n_55100_56840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2089 n_53580_73640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2090 n_55100_70840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2091 n_53580_70840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2092 n_55100_73640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2093 n_58520_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2094 n_61560_73640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2095 n_56620_73640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2096 n_66880_73640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2097 n_58140_79240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2098 n_74100_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2099 n_75240_65240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2100 n_55480_48440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2101 n_40280_73640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2102 n_68780_70840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2103 n_53580_65240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2104 n_53580_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2105 n_54720_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2106 n_48640_79240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2107 n_60040_76440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2108 n_60040_79240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2109 n_63080_79240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2110 n_67260_70840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2111 n_49020_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2112 n_46360_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2113 n_44840_70840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2114 n_44840_76440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2115 n_41800_70840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2116 n_40660_79240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2117 n_43700_79240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2118 n_63080_76440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2119 n_80560_76440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2120 n_54720_84840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2121 n_47120_82040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2122 n_53580_82040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2123 n_40280_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2124 n_52820_79240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2125 n_46740_84840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2126 n_61940_84840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2127 n_49400_84840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2128 n_50920_87640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2129 n_59660_84840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2130 n_55100_82040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2131 n_42940_54040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2132 n_41800_65240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2133 n_43320_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2134 n_43320_76440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2135 n_44080_82040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2136 n_65360_59640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2137 n_65360_56840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2138 n_63080_54040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2139 n_68780_56840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2140 n_59280_87640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2141 n_51680_84840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2142 n_74860_87640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2143 n_54340_87640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2144 n_58520_84840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2145 n_73340_87640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2146 n_56240_76440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2147 n_65360_65240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2148 n_63460_62440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2149 n_63460_59640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2150 n_63460_56840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2151 n_60040_54040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2152 n_67260_56840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2153 n_71820_59640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2154 n_70300_65240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2155 n_71820_65240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2156 n_71820_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2157 n_73720_65240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2158 n_70300_70840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2159 n_70300_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2160 n_67260_76440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2161 n_68780_76440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2162 n_56620_84840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2163 n_87020_59640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2164 n_83220_62440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2165 n_83220_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2166 n_84740_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2167 n_83600_70840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2168 n_85500_70840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2169 n_85880_68040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2170 n_85880_73640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2171 n_83600_76440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2172 n_85500_76440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2173 n_85500_79240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2174 n_83600_79240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2175 n_85500_82040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2176 n_69920_82040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2177 n_68780_82040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2178 n_72200_82040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2179 n_43320_65240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2180 n_40280_62440 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2181 n_60040_56840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2182 n_60040_59640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I2183 n_93480_62440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2184 n_91200_70840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2185 n_91960_87640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2186 n_87020_87640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2187 n_93480_56840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2188 n_93480_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2189 n_93480_76440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2190 n_65740_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2191 n_63840_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2192 n_79040_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2193 n_93480_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2194 n_93480_54040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2195 n_92340_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2196 n_41800_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2197 n_50920_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2198 n_70300_40040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2199 n_87020_40040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2200 n_88160_40040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2201 n_90440_40040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2202 n_93480_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2203 n_80560_40040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2204 n_40280_40040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2205 n_60040_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2206 n_72200_40040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2207 n_82080_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2208 n_43320_59640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2209 n_42180_73640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2210 n_45600_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2211 n_40660_65240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2212 n_47500_40040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2213 n_41800_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2214 n_47500_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2215 n_52060_73640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2216 n_46740_59640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2217 n_80180_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2218 n_71820_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2219 n_56620_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2220 n_41420_40040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2221 n_80180_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2222 n_88920_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2223 n_83600_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2224 n_83600_40040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2225 n_87020_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2226 n_68400_40040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2227 n_51680_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2228 n_48260_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2229 n_85120_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2230 n_92340_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2231 n_90440_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2232 n_78280_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2233 n_64980_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2234 n_64600_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2235 n_90440_76440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2236 n_92340_65240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2237 n_88920_56840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2238 n_85120_84840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2239 n_87400_84840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2240 n_87400_73640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2241 n_91580_62440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2242 n_73340_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2243 n_71820_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2244 n_73340_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2245 n_68780_79240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2246 n_83220_54040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2247 n_91200_54040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2248 n_90820_65240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2249 n_88920_70840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2250 n_87400_65240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2251 n_87400_70840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2252 n_92720_82040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2253 n_92340_76440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2254 n_88920_82040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2255 n_83600_84840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2256 n_83600_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2257 n_80560_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2258 n_85500_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2259 n_84740_54040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2260 n_87400_56840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2261 n_88920_65240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2262 n_88920_76440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2263 n_80560_54040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2264 n_77900_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2265 n_82080_54040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2266 n_80560_56840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2267 n_82080_56840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2268 n_83600_56840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2269 n_76380_54040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2270 n_80560_65240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2271 n_77900_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2272 n_76000_70840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2273 n_79040_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2274 n_74860_70840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2275 n_88920_79240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2276 n_70300_87640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2277 n_70300_84840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2278 n_72200_84840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2279 n_82080_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2280 n_85500_56840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2281 n_86260_54040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2282 n_87400_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2283 n_82080_59640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2284 n_85500_59640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2285 n_84740_65240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2286 n_82080_65240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2287 n_82080_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2288 n_85880_65240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2289 n_87400_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2290 n_80560_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2291 n_77140_70840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2292 n_80560_73640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2293 n_81700_76440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2294 n_79040_70840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2295 n_78660_76440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2296 n_78660_79240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2297 n_76760_76440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2298 n_72200_76440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2299 n_76760_79240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2300 n_80560_79240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2301 n_71820_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2302 n_71820_54040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2303 n_53580_54040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2304 n_68020_54040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2305 n_68780_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2306 n_59280_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2307 n_61940_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2308 n_47880_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2309 n_50920_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2310 n_70300_54040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2311 n_61560_54040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2312 n_66120_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2313 n_76380_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2314 n_76760_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2315 n_90820_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2316 n_90820_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2317 n_85500_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2318 n_50160_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2319 n_51680_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2320 n_46360_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2321 n_48260_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2322 n_70300_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2323 n_87400_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2324 n_85500_40040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2325 n_50540_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2326 n_49400_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2327 n_46740_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2328 n_43320_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2329 n_61560_40040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2330 n_57380_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2331 n_68020_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2332 n_68780_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2333 n_85500_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2334 n_88920_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2335 n_73720_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2336 n_43320_40040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2337 n_58520_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2338 n_73720_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2339 n_76760_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2340 n_74860_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2341 n_80560_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2342 n_53200_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2343 n_55100_62440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2344 n_44080_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2345 n_46740_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2346 n_43320_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2347 n_45220_54040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2348 n_48640_59640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2349 n_48260_65240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2350 n_44840_73640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2351 n_50160_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2352 n_51680_76440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2353 n_40280_59640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2354 n_72200_56840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2355 n_49400_65240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2356 n_56620_65240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2357 n_61560_62440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2358 n_61560_65240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2359 n_60420_65240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2360 n_73720_62440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2361 n_66880_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2362 n_76380_62440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2363 n_63080_82040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2364 n_77520_62440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2365 n_72200_62440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2366 n_73340_59640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2367 n_55100_56840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2368 n_53580_73640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2369 n_50920_73640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2370 n_55860_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2371 n_46740_73640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2372 n_40660_76440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2373 n_40660_70840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2374 n_50920_79240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2375 n_46360_79240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2376 n_58520_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2377 n_70300_73640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2378 n_63460_70840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2379 n_65360_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2380 n_68780_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2381 n_75240_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2382 n_75240_65240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2383 n_72960_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2384 n_55480_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2385 n_40280_73640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2386 n_68780_70840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2387 n_46740_70840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2388 n_48260_76440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2389 n_47500_79240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2390 n_45600_84840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2391 n_58520_70840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2392 n_49400_79240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2393 n_60420_70840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2394 n_76760_73640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2395 n_70300_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2396 n_49020_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2397 n_40660_79240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2398 n_40280_82040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2399 n_43700_79240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2400 n_44080_84840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2401 n_40280_87640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2402 n_80560_76440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2403 n_54720_84840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2404 n_47120_82040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2405 n_50160_84840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2406 n_65740_73640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2407 n_70300_76440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2408 n_47500_56840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2409 n_40280_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2410 n_52820_79240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2411 n_43320_87640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2412 n_46740_84840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2413 n_61940_84840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2414 n_52440_87640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2415 n_49400_87640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2416 n_64220_82040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2417 n_58140_87640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2418 n_42940_54040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2419 n_41800_65240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2420 n_65360_59640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2421 n_65360_56840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2422 n_59280_87640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2423 n_60800_84840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2424 n_60800_87640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2425 n_54340_76440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2426 n_54340_87640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2427 n_65740_82040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2428 n_53580_87640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2429 n_58520_84840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2430 n_64600_84840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2431 n_63460_87640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2432 n_65360_65240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2433 n_63460_62440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2434 n_60040_54040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2435 n_66880_59640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2436 n_71820_59640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2437 n_70300_65240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2438 n_71820_65240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2439 n_71820_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2440 n_73720_65240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2441 n_70300_70840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2442 n_70300_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2443 n_67260_76440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2444 n_65740_79240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2445 n_64600_79240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2446 n_57380_82040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2447 n_55100_79240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2448 n_87400_62440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2449 n_88920_62440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2450 n_87020_59640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2451 n_88160_59640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2452 n_85880_62440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2453 n_83220_65240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2454 n_83220_62440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2455 n_83220_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2456 n_84740_68040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2457 n_83600_70840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2458 n_85500_70840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2459 n_84740_73640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2460 n_83600_76440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2461 n_85500_76440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2462 n_87400_82040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2463 n_71060_82040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2464 n_40280_62440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2465 n_44460_56840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2466 n_60040_56840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I2467 n_92340_54040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2468 n_90820_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2469 n_93480_79240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2470 n_93480_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2471 n_93100_84840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2472 n_83600_87640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2473 n_84740_87640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2474 n_65740_40040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2475 n_65740_45640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2476 n_61940_48440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2477 n_40280_54040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2478 n_44080_54040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2479 n_40660_56840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2480 n_93480_48440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2481 n_41800_42840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2482 n_48640_40040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2483 n_50920_48440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2484 n_63840_40040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2485 n_91580_40040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2486 n_52440_40040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2487 n_80560_40040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2488 n_40280_40040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2489 n_60040_45640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2490 n_72200_40040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2491 n_79040_40040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2492 n_77140_40040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2493 n_40660_45640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2494 n_40660_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2495 n_50160_59640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2496 n_42180_73640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2497 n_44460_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2498 n_43320_62440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2499 n_44460_62440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2500 n_46740_65240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2501 n_52060_73640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2502 n_51300_59640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2503 n_44840_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2504 n_45220_48440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2505 n_74860_40040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2506 n_76760_42840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2507 n_71820_42840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2508 n_56620_45640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2509 n_41420_40040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2510 n_80180_42840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2511 n_51680_42840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2512 n_92720_40040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2513 n_63460_42840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2514 n_51680_48440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2515 n_47880_42840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2516 n_48260_45640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2517 n_90440_48440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2518 n_41420_54040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2519 n_49020_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2520 n_47880_54040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2521 n_60040_48440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2522 n_64600_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2523 n_63080_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2524 n_81700_87640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2525 n_80180_87640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2526 n_90820_84840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2527 n_92340_65240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2528 n_91580_79240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2529 n_88540_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2530 n_89300_54040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2531 n_68780_79240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2532 n_88920_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2533 n_87400_65240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2534 n_92340_76440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2535 n_88920_65240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2536 n_89300_84840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2537 n_80560_84840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2538 n_81700_82040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2539 n_80560_65240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2540 n_77900_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2541 n_76000_70840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2542 n_79040_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2543 n_74860_70840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2544 n_75240_76440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2545 n_73720_79240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2546 n_70300_79240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2547 n_67260_84840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2548 n_88920_79240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2549 n_65740_84840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2550 n_62320_82040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2551 n_65360_87640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2552 n_68780_87640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2553 n_68780_84840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2554 n_70300_84840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2555 n_73720_82040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2556 n_72200_84840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2557 n_86260_54040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2558 n_87400_48440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2559 n_85500_59640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2560 n_84740_65240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2561 n_82080_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2562 n_85880_65240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2563 n_87400_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2564 n_80560_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2565 n_77140_70840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2566 n_78660_76440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2567 n_78660_79240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2568 n_76760_76440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2569 n_76760_79240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2570 n_80180_82040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2571 n_76760_84840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2572 n_76380_87640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2573 n_67260_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2574 n_71820_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2575 n_71820_54040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2576 n_53580_54040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2577 n_68020_54040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2578 n_68780_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2579 n_59280_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2580 n_49780_54040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2581 n_47880_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2582 n_52060_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2583 n_70300_54040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2584 n_61560_54040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2585 n_87400_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2586 n_49400_48440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2587 n_51680_45640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2588 n_53200_48440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2589 n_65360_42840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2590 n_92720_42840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2591 n_50540_42840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2592 n_82080_42840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2593 n_43320_40040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2594 n_53200_45640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2595 n_73720_45640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2596 n_76760_45640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2597 n_73340_40040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2598 n_44080_48440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2599 n_43320_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2600 n_57000_54040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2601 n_52060_54040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2602 n_48260_65240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2603 n_59660_62440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2604 n_44840_73640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2605 n_50160_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2606 n_51680_76440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2607 n_72200_56840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2608 n_53580_59640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2609 n_53580_62440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2610 n_52060_65240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2611 n_49400_65240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2612 n_56620_65240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2613 n_61560_62440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2614 n_61560_65240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2615 n_60420_65240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2616 n_73720_62440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2617 n_66880_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2618 n_76380_62440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2619 n_63080_82040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2620 n_72200_62440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2621 n_73340_59640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2622 n_55100_56840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2623 n_55100_70840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2624 n_53580_70840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2625 n_50920_70840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2626 n_50920_73640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2627 n_55860_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2628 n_46740_73640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2629 n_40660_76440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2630 n_40660_70840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2631 n_50920_79240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2632 n_46360_79240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2633 n_58520_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2634 n_70300_73640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2635 n_63460_70840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2636 n_65360_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2637 n_68780_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2638 n_75240_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2639 n_75240_65240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2640 n_72960_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2641 n_68780_70840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2642 n_53580_65240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2643 n_53580_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2644 n_49400_70840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2645 n_46740_70840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2646 n_48260_76440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2647 n_47500_79240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2648 n_45600_84840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2649 n_58520_70840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2650 n_49400_79240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2651 n_60420_70840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2652 n_76760_73640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2653 n_63080_79240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2654 n_61560_79240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2655 n_65740_76440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2656 n_58140_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2657 n_40660_79240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2658 n_40280_82040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2659 n_43700_79240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2660 n_40280_87640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2661 n_57380_76440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2662 n_63080_76440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2663 n_80560_76440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2664 n_70300_76440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2665 n_47500_56840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2666 n_52820_79240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2667 n_44080_59640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2668 n_42940_82040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2669 n_42940_84840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2670 n_40280_84840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2671 n_43320_87640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2672 n_52440_87640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2673 n_58140_87640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2674 n_65360_62440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2675 n_65360_54040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2676 n_65360_56840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2677 n_63080_54040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2678 n_45220_87640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2679 n_59280_87640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2680 n_51680_84840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2681 n_60800_84840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2682 n_60800_87640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2683 n_54340_76440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2684 n_54340_87640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2685 n_67260_82040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2686 n_65740_82040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2687 n_53580_87640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2688 n_58520_84840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2689 n_64600_84840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2690 n_63460_87640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2691 n_65360_65240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2692 n_63460_62440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2693 n_71820_59640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2694 n_70300_65240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2695 n_71820_65240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2696 n_71820_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2697 n_73720_65240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2698 n_70300_70840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2699 n_70300_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2700 n_67260_76440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2701 n_65740_79240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2702 n_53960_79240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2703 n_55100_79240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2704 n_58520_82040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2705 n_59660_82040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2706 n_87400_62440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2707 n_87020_59640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2708 n_88160_59640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2709 n_83220_65240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2710 n_84740_62440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2711 n_83220_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2712 n_84740_68040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2713 n_83600_70840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2714 n_85500_70840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2715 n_84740_73640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2716 n_85880_73640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2717 n_83600_76440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2718 n_85500_76440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2719 n_87400_82040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2720 n_71060_82040 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2721 n_60040_59640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I2722 n_93480_62440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2723 n_91200_70840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2724 n_93480_79240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2725 n_87020_87640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2726 n_93480_56840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2727 n_90440_62440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2728 n_93480_68040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2729 n_93100_84840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2730 n_56240_48440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2731 n_61940_48440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2732 n_44080_54040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2733 n_40660_56840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2734 n_93480_48440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2735 n_92340_48440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2736 n_48640_40040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2737 n_50920_48440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2738 n_91580_40040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2739 n_87020_40040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2740 n_88160_40040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2741 n_52440_40040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2742 n_40660_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2743 n_42940_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2744 n_90440_40040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2745 n_93480_45640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2746 n_80560_40040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2747 n_40280_48440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2748 n_60040_45640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2749 n_72200_40040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2750 n_82080_48440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2751 n_77140_40040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2752 n_55100_40040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2753 n_40660_51240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2754 n_42180_73640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2755 n_44460_68040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2756 n_46740_65240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2757 n_52060_73640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2758 n_44840_51240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2759 n_54720_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2760 n_74860_40040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2761 n_80180_45640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2762 n_71820_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2763 n_56620_45640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2764 n_41420_48440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2765 n_80180_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2766 n_88920_45640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2767 n_83600_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2768 n_44840_45640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2769 n_43700_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2770 n_51680_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2771 n_83600_40040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2772 n_87020_45640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2773 n_92720_40040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2774 n_51680_48440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2775 n_47880_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2776 n_85120_48440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2777 n_90440_48440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2778 n_41420_54040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2779 n_49020_51240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2780 n_60040_48440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2781 n_55100_54040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2782 n_90820_84840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2783 n_92340_65240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2784 n_90820_59640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2785 n_88920_56840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2786 n_85120_84840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2787 n_91580_79240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2788 n_87400_73640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2789 n_91580_62440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2790 n_87780_54040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2791 n_88920_51240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2792 n_83220_54040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2793 n_91200_54040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2794 n_90820_65240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2795 n_87400_70840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2796 n_92720_82040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2797 n_87780_87640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2798 n_88920_82040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2799 n_83600_84840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2800 n_83600_51240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2801 n_80560_51240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2802 n_84740_54040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2803 n_87400_56840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2804 n_77520_54040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2805 n_87400_79240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2806 n_92720_59640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2807 n_88920_65240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2808 n_89300_73640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2809 n_92340_73640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2810 n_89300_84840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2811 n_81700_82040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2812 n_79040_87640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2813 n_79040_54040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2814 n_80560_54040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2815 n_82080_54040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2816 n_80180_59640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2817 n_79040_68040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2818 n_75240_73640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2819 n_74860_70840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2820 n_75240_76440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2821 n_71820_79240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2822 n_88920_79240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2823 n_67260_87640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2824 n_65360_87640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2825 n_70300_84840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2826 n_73720_82040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2827 n_72200_84840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2828 n_85500_56840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2829 n_82080_59640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2830 n_82080_65240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2831 n_85880_65240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2832 n_77140_70840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2833 n_80560_73640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2834 n_79040_70840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2835 n_72200_76440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2836 n_80180_82040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2837 n_76760_84840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2838 n_76380_87640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2839 n_74860_84840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2840 n_68020_54040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2841 n_61940_51240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2842 n_50920_51240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2843 n_52060_51240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2844 n_87400_51240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2845 n_83600_48440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2846 n_51680_45640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2847 n_53200_48440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2848 n_92720_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2849 n_90440_45640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2850 n_85500_40040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2851 n_50540_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2852 n_45220_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2853 n_46740_45640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2854 n_85500_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2855 n_88920_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2856 n_82080_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2857 n_42940_48440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2858 n_53200_45640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2859 n_73720_45640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2860 n_82080_45640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2861 n_73340_40040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2862 n_53200_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2863 n_43320_51240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2864 n_58900_48440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2865 n_52060_54040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2866 n_66880_68040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2867 n_77520_62440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2868 n_55100_70840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2869 n_53580_70840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2870 n_50920_70840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2871 n_50920_73640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2872 n_49400_73640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2873 n_55860_68040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2874 n_46360_76440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2875 n_48260_73640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2876 n_49780_76440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2877 n_50920_79240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2878 n_58520_68040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2879 n_56620_73640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2880 n_66880_73640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2881 n_74100_68040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2882 n_75240_65240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2883 n_68780_70840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2884 n_53580_65240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2885 n_53580_68040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2886 n_49400_70840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2887 n_46740_70840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2888 n_48260_76440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2889 n_47500_79240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2890 n_58520_70840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2891 n_60420_70840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2892 n_63080_73640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2893 n_63080_79240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2894 n_61560_79240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2895 n_65740_76440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2896 n_67260_70840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2897 n_58140_51240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2898 n_70300_48440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2899 n_57380_76440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2900 n_63080_76440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2901 n_80560_76440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2902 n_65740_73640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2903 n_52440_87640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2904 n_49400_87640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2905 n_64220_82040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2906 n_58140_87640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2907 n_42940_54040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2908 n_46740_51240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2909 n_74860_87640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2910 n_54340_87640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2911 n_67260_82040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2912 n_53580_87640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2913 n_73340_87640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2914 n_57000_87640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2915 n_73720_65240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2916 n_70300_68040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2917 n_59660_82040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2918 n_56240_82040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2919 n_88920_62440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2920 n_87020_59640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2921 n_85880_62440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2922 n_84740_62440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2923 n_83220_62440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2924 n_83600_70840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2925 n_83220_73640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2926 n_85880_73640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2927 n_68780_82040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2928 n_71060_82040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2929 n_43320_65240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2930 n_44460_56840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I2931 n_91200_70840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2932 n_93480_79240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2933 n_93100_87640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2934 n_93480_56840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2935 n_90440_62440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2936 n_93480_73640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2937 n_84740_87640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2938 n_65740_45640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2939 n_61940_48440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2940 n_40280_54040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2941 n_44080_54040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2942 n_93480_54040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2943 n_92340_48440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2944 n_41800_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2945 n_48640_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2946 n_63840_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2947 n_70300_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2948 n_91580_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2949 n_87020_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2950 n_88160_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2951 n_52440_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2952 n_40660_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2953 n_42940_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2954 n_56620_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2955 n_67260_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2956 n_40280_48440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2957 n_72200_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2958 n_82080_48440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2959 n_55100_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2960 n_40660_45640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2961 n_50160_59640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2962 n_43320_62440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2963 n_44460_62440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2964 n_51300_59640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2965 n_45220_48440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2966 n_54720_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2967 n_80180_45640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2968 n_71820_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2969 n_41420_48440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2970 n_66880_45640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2971 n_57760_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2972 n_44840_45640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2973 n_43700_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2974 n_51680_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2975 n_83600_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2976 n_87020_45640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2977 n_92720_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2978 n_68400_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2979 n_63460_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2980 n_47880_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2981 n_48260_45640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2982 n_85120_48440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2983 n_92340_51240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2984 n_49020_51240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2985 n_47880_54040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2986 n_60040_48440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2987 n_64600_51240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2988 n_81700_87640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2989 n_90440_73640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2990 n_90820_59640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2991 n_88920_56840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2992 n_90060_87640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2993 n_91580_79240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2994 n_87400_73640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2995 n_87780_54040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2996 n_88920_51240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2997 n_83220_54040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2998 n_91200_54040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I2999 n_87400_70840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3000 n_92720_82040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3001 n_87780_87640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3002 n_88920_82040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3003 n_83600_84840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3004 n_82080_84840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3005 n_85880_87640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3006 n_83600_51240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3007 n_80560_51240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3008 n_84740_54040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3009 n_87400_56840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3010 n_77520_54040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3011 n_87400_79240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3012 n_92720_59640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3013 n_92340_73640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3014 n_79040_87640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3015 n_79040_54040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3016 n_80560_54040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3017 n_82080_54040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3018 n_82080_56840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3019 n_78660_56840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3020 n_76760_65240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3021 n_78660_65240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3022 n_80560_65240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3023 n_73720_70840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3024 n_71820_79240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3025 n_65740_84840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3026 n_62320_82040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3027 n_70300_87640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3028 n_70300_84840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3029 n_73720_82040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3030 n_85500_56840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3031 n_85500_59640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3032 n_84740_65240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3033 n_82080_68040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3034 n_82080_70840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3035 n_81700_73640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3036 n_80560_73640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3037 n_78660_73640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3038 n_78660_76440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3039 n_78660_79240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3040 n_72200_76440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3041 n_78280_82040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3042 n_76760_79240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3043 n_80180_82040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3044 n_74860_82040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3045 n_76760_82040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3046 n_68780_51240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3047 n_61940_51240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3048 n_49780_54040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3049 n_50920_51240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3050 n_90820_51240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3051 n_83600_48440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3052 n_49400_48440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3053 n_51680_45640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3054 n_65360_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3055 n_70300_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3056 n_92720_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3057 n_90440_45640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3058 n_85500_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3059 n_50540_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3060 n_45220_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3061 n_46740_45640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3062 n_61560_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3063 n_68020_48440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3064 n_42940_48440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3065 n_73720_45640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3066 n_82080_45640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3067 n_53200_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3068 n_44080_48440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3069 n_58900_48440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3070 n_57000_54040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3071 n_48260_65240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3072 n_49780_62440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3073 n_44840_73640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3074 n_50160_68040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3075 n_51680_76440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3076 n_53580_59640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3077 n_53580_62440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3078 n_52060_65240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3079 n_49400_65240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3080 n_56620_65240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3081 n_58520_65240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3082 n_59660_68040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3083 n_60800_68040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3084 n_63460_68040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3085 n_60040_73640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3086 n_63080_65240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3087 n_61940_68040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3088 n_59660_70840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3089 n_55100_56840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3090 n_69160_62440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3091 n_49400_73640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3092 n_46740_73640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3093 n_46360_76440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3094 n_40660_76440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3095 n_48260_73640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3096 n_40660_70840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3097 n_49780_76440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3098 n_46360_79240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3099 n_58520_68040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3100 n_61560_73640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3101 n_58520_73640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3102 n_70300_73640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3103 n_58140_79240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3104 n_63460_70840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3105 n_65360_68040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3106 n_68780_68040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3107 n_68020_62440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3108 n_45600_84840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3109 n_49400_79240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3110 n_63080_73640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3111 n_71820_73640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3112 n_56620_79240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3113 n_60040_79240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3114 n_63080_79240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3115 n_52060_82040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3116 n_40660_79240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3117 n_40280_82040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3118 n_43700_79240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3119 n_40280_87640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3120 n_57380_76440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3121 n_63080_76440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3122 n_80560_76440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3123 n_50920_82040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3124 n_49400_82040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3125 n_54720_84840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3126 n_53580_82040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3127 n_47500_56840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3128 n_52820_79240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3129 n_44080_59640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3130 n_42940_82040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3131 n_42940_84840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3132 n_40280_84840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3133 n_43320_87640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3134 n_46740_84840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3135 n_61940_84840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3136 n_49400_84840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3137 n_49400_87640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3138 n_64220_82040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3139 n_55100_82040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3140 n_45220_87640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3141 n_59280_87640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3142 n_51680_84840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3143 n_60800_84840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3144 n_61180_82040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3145 n_54340_76440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3146 n_67260_82040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3147 n_73340_87640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3148 n_71820_59640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3149 n_70300_65240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3150 n_68400_65240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3151 n_71820_65240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3152 n_71820_68040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3153 n_70300_70840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3154 n_71820_70840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3155 n_67260_76440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3156 n_68780_76440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3157 n_65740_79240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3158 n_53960_79240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3159 n_55100_79240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3160 n_59660_82040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3161 n_83600_70840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3162 n_83220_73640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3163 n_85880_73640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3164 n_81700_79240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3165 n_43320_65240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3166 n_44460_56840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I3167 n_92340_54040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3168 n_93480_62440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3169 n_93480_79240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3170 n_91960_87640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3171 n_90440_62440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3172 n_65740_40040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3173 n_54720_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3174 n_61940_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3175 n_44080_54040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3176 n_40660_56840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3177 n_63840_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3178 n_79040_42840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3179 n_92340_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3180 n_48640_40040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3181 n_50920_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3182 n_63840_40040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3183 n_91580_40040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3184 n_87020_40040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3185 n_52440_40040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3186 n_42940_42840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3187 n_67260_40040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3188 n_90440_40040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3189 n_40280_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3190 n_60040_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3191 n_72200_40040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3192 n_82080_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3193 n_44460_68040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3194 n_43320_62440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3195 n_44460_62440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3196 n_46740_65240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3197 n_80180_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3198 n_71820_42840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3199 n_56620_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3200 n_41420_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3201 n_83600_42840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3202 n_66880_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3203 n_44840_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3204 n_51680_42840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3205 n_87020_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3206 n_92720_40040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3207 n_63460_42840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3208 n_51680_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3209 n_47880_42840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3210 n_85120_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3211 n_78280_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3212 n_64980_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3213 n_41420_54040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3214 n_49020_51240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3215 n_60040_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3216 n_54720_51240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3217 n_63080_51240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3218 n_90820_59640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3219 n_87400_84840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3220 n_91580_79240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3221 n_91580_62440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3222 n_89300_54040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3223 n_88920_51240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3224 n_83220_54040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3225 n_91200_54040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3226 n_92340_56840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3227 n_92720_82040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3228 n_88920_82040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3229 n_83600_84840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3230 n_82080_84840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3231 n_88920_87640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3232 n_85880_87640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3233 n_83600_51240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3234 n_80560_51240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3235 n_84740_54040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3236 n_87400_56840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3237 n_90820_56840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3238 n_77520_54040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3239 n_87400_79240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3240 n_92720_59640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3241 n_79040_54040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3242 n_80560_54040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3243 n_82080_54040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3244 n_80560_56840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3245 n_80180_59640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3246 n_83600_56840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3247 n_76380_54040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3248 n_76760_56840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3249 n_71820_79240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3250 n_70300_87640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3251 n_70300_84840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3252 n_73720_82040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3253 n_85500_56840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3254 n_87400_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3255 n_85500_59640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3256 n_87400_68040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3257 n_80560_68040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3258 n_81700_73640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3259 n_80560_70840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3260 n_80560_73640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3261 n_81700_76440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3262 n_78660_73640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3263 n_78660_76440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3264 n_78660_79240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3265 n_72200_76440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3266 n_78280_82040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3267 n_76760_79240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3268 n_80560_79240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3269 n_80180_82040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3270 n_76760_84840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3271 n_76380_87640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3272 n_74860_84840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3273 n_74860_82040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3274 n_76760_82040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3275 n_67260_51240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3276 n_70300_51240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3277 n_61940_51240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3278 n_50920_51240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3279 n_52060_51240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3280 n_66120_51240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3281 n_79040_51240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3282 n_83600_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3283 n_51680_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3284 n_53200_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3285 n_65360_42840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3286 n_92720_42840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3287 n_90440_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3288 n_50540_42840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3289 n_46740_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3290 n_68020_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3291 n_85500_42840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3292 n_42940_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3293 n_53200_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3294 n_73720_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3295 n_82080_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3296 n_58900_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3297 n_57000_54040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3298 n_52060_54040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3299 n_49780_62440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3300 n_59660_62440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3301 n_44840_73640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3302 n_50920_68040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3303 n_50160_68040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3304 n_51680_76440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3305 n_72200_56840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3306 n_61560_62440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3307 n_75240_59640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3308 n_77520_62440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3309 n_72200_62440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3310 n_55100_56840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3311 n_49400_73640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3312 n_46740_73640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3313 n_40660_76440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3314 n_48260_73640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3315 n_40660_70840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3316 n_49780_76440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3317 n_46360_79240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3318 n_61560_73640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3319 n_58140_79240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3320 n_55480_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3321 n_53580_65240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3322 n_53580_68040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3323 n_54720_68040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3324 n_46740_70840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3325 n_48260_76440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3326 n_47500_79240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3327 n_45600_84840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3328 n_58520_70840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3329 n_49400_79240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3330 n_60420_70840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3331 n_63080_73640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3332 n_56620_79240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3333 n_60040_79240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3334 n_63080_79240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3335 n_65740_76440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3336 n_58140_51240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3337 n_70300_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3338 n_40660_79240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3339 n_40280_82040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3340 n_43700_79240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3341 n_44080_84840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3342 n_57380_76440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3343 n_63080_76440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3344 n_50920_82040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3345 n_50160_84840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3346 n_65740_73640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3347 n_47500_56840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3348 n_44080_59640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3349 n_42940_82040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3350 n_45220_82040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3351 n_40280_84840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3352 n_41420_87640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3353 n_46740_87640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3354 n_43320_87640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3355 n_46740_84840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3356 n_52440_87640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3357 n_49400_87640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3358 n_64220_82040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3359 n_58140_87640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3360 n_46740_51240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3361 n_65360_62440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3362 n_65360_54040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3363 n_65360_56840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3364 n_68780_56840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3365 n_59280_87640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3366 n_60800_84840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3367 n_61180_82040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3368 n_74860_87640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3369 n_54340_76440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3370 n_54340_87640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3371 n_67260_82040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3372 n_53580_87640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3373 n_57000_87640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3374 n_65360_65240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3375 n_63460_62440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3376 n_63460_59640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3377 n_63460_56840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3378 n_68780_59640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3379 n_67260_56840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3380 n_66880_59640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3381 n_70300_59640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3382 n_70300_56840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3383 n_71820_59640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3384 n_67260_76440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3385 n_68780_76440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3386 n_65740_79240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3387 n_64600_79240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3388 n_64600_76440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3389 n_58520_82040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3390 n_59660_82040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3391 n_56240_82040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3392 n_88920_62440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3393 n_87020_59640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3394 n_84740_68040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3395 n_85880_73640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3396 n_85500_82040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3397 n_68780_82040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I3398 n_91200_70840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3399 n_93100_87640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3400 n_93480_56840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3401 n_90440_62440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3402 n_93480_68040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3403 n_93480_73640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3404 n_93100_84840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3405 n_84740_87640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3406 n_54720_48440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3407 n_56240_48440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3408 n_65740_45640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3409 n_79040_42840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3410 n_93480_48440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3411 n_93480_54040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3412 n_63840_40040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3413 n_87020_40040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3414 n_42940_42840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3415 n_67260_40040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3416 n_90440_40040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3417 n_93480_45640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3418 n_46360_40040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3419 n_82080_48440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3420 n_44460_68040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3421 n_45600_68040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3422 n_40660_65240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3423 n_41800_68040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3424 n_47500_68040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3425 n_46740_65240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3426 n_80180_45640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3427 n_49400_40040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3428 n_88920_45640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3429 n_83600_42840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3430 n_66880_45640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3431 n_44840_45640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3432 n_87020_45640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3433 n_63460_42840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3434 n_92340_51240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3435 n_90440_48440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3436 n_78280_48440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3437 n_64600_51240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3438 n_55100_54040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3439 n_54720_51240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3440 n_81700_87640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3441 n_90820_84840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3442 n_90440_73640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3443 n_92340_65240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3444 n_90820_59640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3445 n_88920_56840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3446 n_90060_87640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3447 n_87400_73640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3448 n_68780_79240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3449 n_83220_54040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3450 n_91200_54040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3451 n_92340_56840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3452 n_90820_65240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3453 n_87400_76440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3454 n_92720_82040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3455 n_92340_76440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3456 n_83600_84840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3457 n_82080_84840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3458 n_88920_87640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3459 n_83600_51240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3460 n_80560_51240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3461 n_84740_54040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3462 n_90820_56840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3463 n_92720_59640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3464 n_91960_68040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3465 n_92340_73640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3466 n_90820_82040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3467 n_79040_87640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3468 n_82080_54040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3469 n_83600_56840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3470 n_76760_56840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3471 n_78280_70840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3472 n_73720_70840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3473 n_67260_84840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3474 n_67260_87640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3475 n_68780_87640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3476 n_68780_84840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3477 n_85500_56840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3478 n_82080_59640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3479 n_84740_65240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3480 n_82080_65240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3481 n_82080_68040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3482 n_85880_65240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3483 n_87400_68040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3484 n_82080_70840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3485 n_80560_68040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3486 n_77140_70840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3487 n_80560_70840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3488 n_81700_76440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3489 n_80180_82040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3490 n_76760_82040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3491 n_70300_51240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3492 n_68020_54040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3493 n_68780_51240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3494 n_79040_51240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3495 n_87400_51240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3496 n_90820_51240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3497 n_65360_42840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3498 n_90440_45640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3499 n_46740_45640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3500 n_68020_48440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3501 n_85500_42840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3502 n_88920_42840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3503 n_51300_40040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3504 n_82080_45640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3505 n_52060_54040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3506 n_61560_65240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3507 n_58520_65240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3508 n_59660_68040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3509 n_60420_65240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3510 n_73720_62440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3511 n_60800_68040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3512 n_63460_68040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3513 n_60040_73640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3514 n_63080_65240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3515 n_76380_62440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3516 n_63080_82040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3517 n_75240_59640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3518 n_73340_59640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3519 n_61940_68040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3520 n_59660_70840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3521 n_46360_76440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3522 n_40660_76440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3523 n_40660_70840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3524 n_58520_68040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3525 n_58520_73640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3526 n_70300_73640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3527 n_66880_73640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3528 n_58140_79240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3529 n_63460_70840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3530 n_65360_70840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3531 n_68780_68040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3532 n_68020_62440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3533 n_53580_65240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3534 n_53580_68040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3535 n_54720_68040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3536 n_48260_76440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3537 n_48640_79240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3538 n_58520_70840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3539 n_60040_76440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3540 n_60420_70840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3541 n_71820_73640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3542 n_56620_79240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3543 n_65740_76440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3544 n_67260_70840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3545 n_46360_68040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3546 n_44840_70840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3547 n_44840_76440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3548 n_40660_79240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3549 n_40280_82040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3550 n_43700_79240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3551 n_44080_84840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3552 n_57380_76440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3553 n_80560_76440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3554 n_53580_82040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3555 n_50160_84840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3556 n_70300_76440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3557 n_47500_56840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3558 n_40280_84840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3559 n_61940_84840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3560 n_63080_84840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3561 n_49400_84840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3562 n_52440_87640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3563 n_58140_87640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3564 n_55100_82040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3565 n_46740_51240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3566 n_43320_68040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3567 n_43320_76440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3568 n_44080_82040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3569 n_63080_54040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3570 n_45220_87640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3571 n_51680_84840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3572 n_74860_87640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3573 n_54340_87640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3574 n_53580_87640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3575 n_58520_84840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3576 n_64600_84840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3577 n_63460_87640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3578 n_63460_59640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3579 n_63460_56840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3580 n_60040_54040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3581 n_70300_65240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3582 n_68400_65240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3583 n_71820_65240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3584 n_71820_68040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3585 n_70300_70840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3586 n_71820_70840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3587 n_58520_82040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3588 n_56240_82040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3589 n_87400_62440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3590 n_87020_59640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3591 n_88160_59640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3592 n_85880_62440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3593 n_83220_65240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3594 n_83220_62440 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3595 n_83220_68040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3596 n_83600_70840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3597 n_83220_73640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3598 n_81700_79240 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3599 n_85500_82040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3600 n_68780_82040 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3601 n_60040_56840 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3602 n_60040_59640 0 PWL(26000ps 0uA 26030ps 0uA 26031ps 30uA 26059ps 30uA 26060ps 0uA)
I3603 n_90820_68040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3604 n_91960_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3605 n_93100_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3606 n_90440_62440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3607 n_93480_76440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3608 n_93100_84840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3609 n_83600_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3610 n_84740_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3611 n_54720_48440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3612 n_79040_42840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3613 n_70300_40040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3614 n_88160_40040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3615 n_42940_42840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3616 n_90440_40040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3617 n_80560_40040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3618 n_60040_45640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3619 n_79040_40040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3620 n_82080_48440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3621 n_77140_40040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3622 n_55100_40040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3623 n_50160_59640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3624 n_45600_68040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3625 n_40660_65240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3626 n_41800_68040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3627 n_47500_68040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3628 n_51300_59640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3629 n_54720_42840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3630 n_74860_40040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3631 n_80180_45640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3632 n_76760_42840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3633 n_56620_45640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3634 n_80180_42840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3635 n_83600_42840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3636 n_44840_45640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3637 n_83600_40040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3638 n_68400_40040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3639 n_78280_48440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3640 n_54720_51240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3641 n_81700_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3642 n_80180_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3643 n_90820_84840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3644 n_90440_76440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3645 n_90820_59640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3646 n_90060_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3647 n_87400_84840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3648 n_88540_68040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3649 n_68780_79240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3650 n_87400_65240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3651 n_88920_82040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3652 n_85880_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3653 n_92720_59640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3654 n_90060_79240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3655 n_90820_82040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3656 n_77900_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3657 n_79040_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3658 n_76760_56840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3659 n_67260_84840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3660 n_71820_79240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3661 n_88920_79240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3662 n_67260_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3663 n_68780_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3664 n_68780_84840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3665 n_70300_84840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3666 n_72200_84840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3667 n_84740_65240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3668 n_82080_68040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3669 n_85880_65240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3670 n_87400_68040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3671 n_82080_70840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3672 n_81700_73640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3673 n_78660_73640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3674 n_78660_76440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3675 n_78660_79240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3676 n_78280_82040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3677 n_76760_79240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3678 n_80560_79240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3679 n_76760_84840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3680 n_76380_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3681 n_74860_84840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3682 n_70300_51240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3683 n_79040_51240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3684 n_70300_42840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3685 n_85500_40040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3686 n_46740_45640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3687 n_85500_42840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3688 n_82080_42840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3689 n_53200_45640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3690 n_76760_45640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3691 n_82080_45640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3692 n_73340_40040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3693 n_53200_42840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3694 n_57000_54040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3695 n_52060_54040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3696 n_48260_65240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3697 n_50920_68040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3698 n_53580_59640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3699 n_53580_62440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3700 n_55100_65240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3701 n_49400_65240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3702 n_56620_65240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3703 n_61560_65240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3704 n_60420_65240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3705 n_73720_62440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3706 n_76380_62440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3707 n_63080_82040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3708 n_75240_59640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3709 n_77520_62440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3710 n_73340_59640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3711 n_40660_76440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3712 n_40660_70840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3713 n_66880_73640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3714 n_58140_79240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3715 n_63460_70840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3716 n_74100_68040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3717 n_65360_70840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3718 n_68780_68040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3719 n_75240_65240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3720 n_68020_62440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3721 n_55480_48440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3722 n_46740_70840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3723 n_47500_79240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3724 n_48640_79240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3725 n_60040_76440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3726 n_56620_79240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3727 n_65740_76440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3728 n_67260_70840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3729 n_46360_68040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3730 n_44840_70840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3731 n_44840_76440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3732 n_40660_79240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3733 n_40280_82040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3734 n_43700_79240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3735 n_40280_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3736 n_57380_76440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3737 n_53580_82040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3738 n_50160_84840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3739 n_70300_76440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3740 n_47500_56840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3741 n_40280_84840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3742 n_41420_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3743 n_43320_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3744 n_61940_84840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3745 n_63080_84840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3746 n_49400_84840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3747 n_52440_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3748 n_59660_84840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3749 n_55100_82040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3750 n_42940_54040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3751 n_43320_68040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3752 n_43320_76440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3753 n_44080_82040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3754 n_63080_54040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3755 n_45220_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3756 n_59280_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3757 n_51680_84840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3758 n_54340_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3759 n_64600_84840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3760 n_56240_76440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3761 n_57000_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3762 n_63460_87640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3763 n_63460_59640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3764 n_63460_56840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3765 n_60040_54040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3766 n_70300_62440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3767 n_58520_82040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3768 n_56240_82040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3769 n_56620_84840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3770 n_84740_62440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3771 n_85500_70840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3772 n_84740_73640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3773 n_85880_68040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3774 n_83600_76440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3775 n_85500_76440 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3776 n_85500_79240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3777 n_83600_82040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3778 n_83600_79240 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3779 n_69920_82040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3780 n_71060_82040 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3781 n_44460_56840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3782 n_60040_56840 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3783 n_60040_59640 0 PWL(28000ps 0uA 28030ps 0uA 28031ps 30uA 28059ps 30uA 28060ps 0uA)
I3784 n_93480_62440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3785 n_93480_79240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3786 n_91960_87640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3787 n_87020_87640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3788 n_93480_56840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3789 n_93480_73640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3790 n_84740_87640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3791 n_65740_40040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3792 n_56240_48440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3793 n_40280_54040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3794 n_44080_54040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3795 n_40660_56840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3796 n_63840_45640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3797 n_92340_48440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3798 n_41800_42840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3799 n_70300_40040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3800 n_88160_40040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3801 n_56620_40040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3802 n_67260_40040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3803 n_93480_45640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3804 n_80560_40040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3805 n_46360_40040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3806 n_72200_40040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3807 n_77140_40040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3808 n_50160_59640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3809 n_44460_68040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3810 n_45600_68040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3811 n_47500_68040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3812 n_46740_65240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3813 n_51300_59640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3814 n_74860_40040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3815 n_71820_42840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3816 n_49400_40040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3817 n_80180_42840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3818 n_88920_45640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3819 n_66880_45640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3820 n_57760_40040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3821 n_83600_40040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3822 n_68400_40040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3823 n_48260_45640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3824 n_85120_48440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3825 n_64980_48440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3826 n_41420_54040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3827 n_49020_51240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3828 n_47880_54040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3829 n_55100_54040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3830 n_63080_51240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3831 n_81700_87640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3832 n_90440_73640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3833 n_88920_56840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3834 n_85120_84840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3835 n_87400_84840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3836 n_91580_79240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3837 n_91580_62440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3838 n_68780_79240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3839 n_90820_65240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3840 n_92340_76440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3841 n_88920_82040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3842 n_82080_84840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3843 n_90820_56840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3844 n_92340_73640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3845 n_79040_87640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3846 n_76380_54040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3847 n_75240_73640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3848 n_74860_70840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3849 n_75240_76440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3850 n_65740_84840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3851 n_62320_82040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3852 n_85500_56840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3853 n_86260_54040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3854 n_82080_59640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3855 n_84740_65240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3856 n_83600_59640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3857 n_82080_65240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3858 n_82080_68040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3859 n_82080_70840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3860 n_81700_73640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3861 n_78660_73640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3862 n_78660_76440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3863 n_78660_79240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3864 n_72200_76440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3865 n_78280_82040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3866 n_76760_79240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3867 n_80560_79240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3868 n_80180_82040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3869 n_76760_84840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3870 n_78660_84840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3871 n_76760_82040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3872 n_60800_51240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3873 n_71820_51240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3874 n_71820_54040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3875 n_53200_51240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3876 n_70300_51240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3877 n_68020_54040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3878 n_56620_51240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3879 n_68780_51240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3880 n_59280_51240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3881 n_61940_51240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3882 n_46360_54040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3883 n_50920_51240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3884 n_52060_51240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3885 n_70300_54040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3886 n_61560_54040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3887 n_66120_51240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3888 n_83600_48440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3889 n_49400_48440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3890 n_70300_42840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3891 n_85500_40040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3892 n_61560_40040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3893 n_68020_48440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3894 n_88920_42840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3895 n_82080_42840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3896 n_51300_40040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3897 n_73720_45640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3898 n_73340_40040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3899 n_58900_48440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3900 n_57000_54040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3901 n_48260_65240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3902 n_50920_68040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3903 n_53580_59640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3904 n_53580_62440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3905 n_55100_65240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3906 n_49400_65240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3907 n_56620_65240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3908 n_61560_65240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3909 n_60420_65240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3910 n_73720_62440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3911 n_66880_68040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3912 n_60800_68040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3913 n_60040_73640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3914 n_76380_62440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3915 n_63080_82040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3916 n_77520_62440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3917 n_59660_70840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3918 n_46360_76440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3919 n_58520_68040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3920 n_61560_73640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3921 n_58140_79240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3922 n_63460_70840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3923 n_65360_70840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3924 n_68780_68040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3925 n_75240_68040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3926 n_75240_65240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3927 n_68020_62440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3928 n_55480_48440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3929 n_68780_70840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3930 n_53580_65240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3931 n_53580_68040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3932 n_54720_68040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3933 n_46740_70840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3934 n_48260_76440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3935 n_47500_79240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3936 n_48640_79240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3937 n_58520_70840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3938 n_60040_76440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3939 n_60420_70840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3940 n_63080_73640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3941 n_60040_79240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3942 n_63080_79240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3943 n_67260_70840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3944 n_68400_73640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3945 n_58140_51240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3946 n_70300_48440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3947 n_46360_68040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3948 n_44840_70840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3949 n_44840_76440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3950 n_41800_70840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3951 n_40660_79240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3952 n_43700_79240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3953 n_67260_79240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3954 n_80560_76440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3955 n_52820_79240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3956 n_61940_84840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3957 n_63080_84840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3958 n_64220_82040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3959 n_50920_87640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3960 n_58140_87640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3961 n_55100_82040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3962 n_61940_87640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3963 n_42940_54040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3964 n_63080_54040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3965 n_68780_56840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3966 n_54340_87640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3967 n_65740_82040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3968 n_53580_87640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3969 n_73340_87640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3970 n_57000_87640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3971 n_63460_59640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3972 n_63460_56840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3973 n_60040_54040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3974 n_68780_59640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3975 n_67260_56840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3976 n_71820_68040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3977 n_73720_65240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3978 n_70300_70840 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3979 n_67260_76440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3980 n_68780_76440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3981 n_53960_79240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3982 n_57380_82040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3983 n_64600_76440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3984 n_55100_79240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3985 n_83220_65240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3986 n_83220_73640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3987 n_84740_73640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3988 n_83600_76440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3989 n_85500_76440 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3990 n_85500_79240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3991 n_83600_82040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3992 n_83600_79240 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3993 n_85500_82040 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3994 n_60040_59640 0 PWL(30000ps 0uA 30030ps 0uA 30031ps 30uA 30059ps 30uA 30060ps 0uA)
I3995 n_93480_62440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I3996 n_90820_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I3997 n_91200_70840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I3998 n_93100_87640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I3999 n_90440_62440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4000 n_93480_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4001 n_93480_76440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4002 n_83600_87640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4003 n_54720_48440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4004 n_65740_45640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4005 n_61940_48440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4006 n_40280_54040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4007 n_44080_54040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4008 n_79040_42840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4009 n_93480_48440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4010 n_93480_54040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4011 n_41800_42840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4012 n_50920_48440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4013 n_63840_40040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4014 n_70300_40040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4015 n_87020_40040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4016 n_88160_40040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4017 n_52440_40040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4018 n_42940_42840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4019 n_67260_40040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4020 n_46360_40040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4021 n_40280_40040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4022 n_60040_45640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4023 n_72200_40040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4024 n_77140_40040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4025 n_55100_40040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4026 n_50160_59640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4027 n_42180_73640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4028 n_44460_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4029 n_45600_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4030 n_43320_62440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4031 n_40660_65240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4032 n_41800_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4033 n_44460_62440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4034 n_47500_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4035 n_46740_65240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4036 n_52060_73640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4037 n_51300_59640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4038 n_54720_42840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4039 n_74860_40040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4040 n_71820_42840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4041 n_56620_45640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4042 n_41420_40040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4043 n_49400_40040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4044 n_66880_45640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4045 n_44840_45640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4046 n_51680_42840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4047 n_83600_40040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4048 n_87020_45640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4049 n_68400_40040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4050 n_63460_42840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4051 n_51680_48440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4052 n_48260_45640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4053 n_92340_51240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4054 n_90440_48440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4055 n_78280_48440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4056 n_49020_51240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4057 n_47880_54040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4058 n_60040_48440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4059 n_64600_51240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4060 n_54720_51240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4061 n_80180_87640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4062 n_90440_76440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4063 n_92340_65240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4064 n_90820_59640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4065 n_90060_87640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4066 n_87400_73640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4067 n_88540_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4068 n_91580_62440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4069 n_68780_79240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4070 n_90820_65240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4071 n_87400_65240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4072 n_87400_76440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4073 n_85880_87640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4074 n_92720_59640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4075 n_91960_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4076 n_90060_79240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4077 n_77900_87640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4078 n_76760_56840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4079 n_78280_70840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4080 n_75240_73640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4081 n_74860_70840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4082 n_73720_70840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4083 n_75240_76440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4084 n_88920_79240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4085 n_65740_84840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4086 n_62320_82040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4087 n_70300_84840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4088 n_72200_84840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4089 n_85500_56840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4090 n_82080_59640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4091 n_83600_59640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4092 n_82080_65240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4093 n_87400_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4094 n_77140_70840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4095 n_80560_73640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4096 n_76760_84840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4097 n_78660_84840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4098 n_74860_84840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4099 n_60800_51240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4100 n_67260_51240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4101 n_71820_51240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4102 n_71820_54040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4103 n_53200_51240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4104 n_56620_51240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4105 n_59280_51240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4106 n_46360_54040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4107 n_50920_51240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4108 n_70300_54040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4109 n_61560_54040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4110 n_79040_51240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4111 n_87400_51240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4112 n_90820_51240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4113 n_49400_48440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4114 n_53200_48440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4115 n_65360_42840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4116 n_70300_42840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4117 n_90440_45640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4118 n_85500_40040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4119 n_50540_42840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4120 n_46740_45640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4121 n_68020_48440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4122 n_51300_40040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4123 n_43320_40040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4124 n_53200_45640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4125 n_73720_45640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4126 n_73340_40040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4127 n_53200_42840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4128 n_58900_48440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4129 n_48260_65240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4130 n_59660_62440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4131 n_50920_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4132 n_53580_59640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4133 n_53580_62440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4134 n_52060_65240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4135 n_49400_65240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4136 n_56620_65240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4137 n_61560_62440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4138 n_61560_65240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4139 n_59660_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4140 n_66880_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4141 n_63080_65240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4142 n_76380_62440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4143 n_75240_62440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4144 n_76380_59640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4145 n_63080_82040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4146 n_77520_62440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4147 n_61940_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4148 n_55100_56840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4149 n_69160_62440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4150 n_55100_70840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4151 n_53580_70840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4152 n_50920_70840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4153 n_50920_73640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4154 n_49400_73640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4155 n_55860_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4156 n_46360_76440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4157 n_49780_76440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4158 n_50920_79240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4159 n_58520_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4160 n_58520_73640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4161 n_70300_73640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4162 n_74100_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4163 n_65360_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4164 n_65360_70840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4165 n_75240_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4166 n_68780_70840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4167 n_53580_65240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4168 n_53580_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4169 n_54720_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4170 n_46740_70840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4171 n_48260_76440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4172 n_47500_79240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4173 n_48640_79240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4174 n_58520_70840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4175 n_60040_76440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4176 n_60420_70840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4177 n_71820_73640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4178 n_56620_79240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4179 n_65740_76440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4180 n_67260_70840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4181 n_68400_73640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4182 n_58140_51240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4183 n_46360_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4184 n_44840_70840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4185 n_44840_76440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4186 n_41800_70840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4187 n_40660_79240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4188 n_43700_79240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4189 n_44080_84840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4190 n_57380_76440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4191 n_63080_76440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4192 n_67260_79240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4193 n_50920_82040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4194 n_50160_84840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4195 n_65740_73640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4196 n_52820_79240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4197 n_44080_59640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4198 n_42940_82040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4199 n_45220_82040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4200 n_40280_84840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4201 n_46740_87640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4202 n_43320_87640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4203 n_46740_84840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4204 n_61940_84840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4205 n_63080_84840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4206 n_52440_87640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4207 n_64220_82040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4208 n_50920_87640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4209 n_58140_87640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4210 n_59660_84840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4211 n_55100_82040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4212 n_61940_87640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4213 n_42940_54040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4214 n_43320_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4215 n_43320_76440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4216 n_41800_82040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4217 n_65360_62440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4218 n_65360_54040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4219 n_65360_56840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4220 n_63080_54040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4221 n_51680_84840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4222 n_60800_84840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4223 n_61180_82040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4224 n_54340_76440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4225 n_65740_82040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4226 n_53580_87640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4227 n_58520_84840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4228 n_73340_87640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4229 n_56240_76440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4230 n_57000_87640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4231 n_65360_65240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4232 n_63460_62440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4233 n_60040_54040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4234 n_66880_59640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4235 n_70300_59640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4236 n_70300_62440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4237 n_70300_56840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4238 n_71820_59640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4239 n_70300_65240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4240 n_71820_65240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4241 n_73720_65240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4242 n_71820_70840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4243 n_65740_79240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4244 n_64600_79240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4245 n_53960_79240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4246 n_57380_82040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4247 n_55100_79240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4248 n_58520_82040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4249 n_56240_82040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4250 n_56620_84840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4251 n_87400_62440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4252 n_87020_59640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4253 n_88160_59640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4254 n_85880_62440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4255 n_84740_62440 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4256 n_83220_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4257 n_84740_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4258 n_83600_70840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4259 n_85500_70840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4260 n_85880_68040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4261 n_85880_73640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4262 n_81700_79240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4263 n_69920_82040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4264 n_68780_82040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4265 n_71060_82040 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4266 n_43320_65240 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4267 n_44460_56840 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4268 n_60040_59640 0 PWL(32000ps 0uA 32030ps 0uA 32031ps 30uA 32059ps 30uA 32060ps 0uA)
I4269 n_90820_68040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4270 n_93480_79240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4271 n_87020_87640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4272 n_93480_56840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4273 n_90440_62440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4274 n_93480_73640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4275 n_93480_76440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4276 n_65740_40040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4277 n_54720_48440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4278 n_65740_45640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4279 n_61940_48440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4280 n_44080_54040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4281 n_40660_56840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4282 n_63840_45640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4283 n_79040_42840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4284 n_93480_54040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4285 n_92340_48440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4286 n_48640_40040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4287 n_50920_48440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4288 n_63840_40040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4289 n_87020_40040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4290 n_88160_40040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4291 n_40660_42840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4292 n_56620_40040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4293 n_67260_40040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4294 n_90440_40040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4295 n_60040_45640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4296 n_72200_40040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4297 n_77140_40040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4298 n_40660_45640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4299 n_42180_73640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4300 n_52060_73640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4301 n_45220_48440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4302 n_74860_40040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4303 n_71820_42840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4304 n_56620_45640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4305 n_83600_42840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4306 n_66880_45640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4307 n_57760_40040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4308 n_43700_42840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4309 n_83600_40040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4310 n_87020_45640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4311 n_63460_42840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4312 n_51680_48440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4313 n_47880_42840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4314 n_85120_48440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4315 n_92340_51240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4316 n_78280_48440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4317 n_64980_48440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4318 n_41420_54040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4319 n_49020_51240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4320 n_60040_48440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4321 n_64600_51240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4322 n_54720_51240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4323 n_63080_51240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4324 n_90440_76440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4325 n_90440_73640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4326 n_90820_59640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4327 n_88920_56840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4328 n_85120_84840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4329 n_91580_79240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4330 n_88540_68040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4331 n_87400_65240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4332 n_92340_76440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4333 n_82080_84840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4334 n_90820_56840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4335 n_77520_54040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4336 n_87400_79240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4337 n_89300_59640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4338 n_89300_73640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4339 n_88920_76440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4340 n_81700_82040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4341 n_79040_87640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4342 n_79040_54040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4343 n_80560_54040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4344 n_80560_56840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4345 n_82080_56840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4346 n_78660_56840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4347 n_76380_54040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4348 n_76760_65240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4349 n_76760_56840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4350 n_76380_68040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4351 n_78280_70840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4352 n_73720_70840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4353 n_67260_84840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4354 n_71820_79240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4355 n_67260_87640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4356 n_68780_87640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4357 n_68780_84840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4358 n_70300_84840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4359 n_73720_82040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4360 n_86260_54040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4361 n_84740_65240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4362 n_82080_68040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4363 n_87400_68040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4364 n_80560_68040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4365 n_79040_70840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4366 n_78660_76440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4367 n_78660_79240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4368 n_72200_76440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4369 n_78280_82040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4370 n_80180_82040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4371 n_74860_84840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4372 n_74860_82040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4373 n_76760_82040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4374 n_67260_51240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4375 n_70300_51240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4376 n_68780_51240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4377 n_61940_51240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4378 n_50920_51240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4379 n_52060_51240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4380 n_66120_51240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4381 n_79040_51240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4382 n_90820_51240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4383 n_83600_48440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4384 n_51680_45640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4385 n_53200_48440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4386 n_65360_42840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4387 n_90440_45640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4388 n_85500_40040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4389 n_45220_42840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4390 n_61560_40040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4391 n_68020_48440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4392 n_85500_42840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4393 n_53200_45640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4394 n_73720_45640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4395 n_73340_40040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4396 n_44080_48440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4397 n_59660_62440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4398 n_55100_65240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4399 n_52060_65240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4400 n_61560_62440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4401 n_59660_68040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4402 n_60420_65240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4403 n_73720_62440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4404 n_60800_68040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4405 n_60040_73640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4406 n_63080_65240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4407 n_75240_62440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4408 n_76380_59640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4409 n_61940_68040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4410 n_59660_70840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4411 n_55100_56840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4412 n_55100_70840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4413 n_53580_70840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4414 n_50920_70840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4415 n_50920_73640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4416 n_49400_73640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4417 n_55860_68040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4418 n_49780_76440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4419 n_50920_79240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4420 n_61560_73640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4421 n_58520_73640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4422 n_70300_73640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4423 n_58140_79240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4424 n_63080_73640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4425 n_71820_73640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4426 n_56620_79240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4427 n_60040_79240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4428 n_63080_79240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4429 n_65740_76440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4430 n_70300_48440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4431 n_57380_76440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4432 n_63080_76440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4433 n_80560_76440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4434 n_65740_73640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4435 n_52440_87640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4436 n_49400_87640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4437 n_64220_82040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4438 n_59660_84840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4439 n_42940_54040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4440 n_44080_82040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4441 n_41800_82040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4442 n_65360_62440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4443 n_65360_54040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4444 n_65360_56840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4445 n_68780_56840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4446 n_60800_84840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4447 n_61180_82040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4448 n_74860_87640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4449 n_54340_76440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4450 n_54340_87640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4451 n_67260_82040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4452 n_58520_84840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4453 n_56240_76440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4454 n_65360_65240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4455 n_63460_62440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4456 n_63460_59640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4457 n_63460_56840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4458 n_68780_59640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4459 n_67260_56840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4460 n_66880_59640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4461 n_70300_59640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4462 n_70300_62440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4463 n_70300_56840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4464 n_71820_59640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4465 n_70300_65240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4466 n_71820_65240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4467 n_71820_68040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4468 n_70300_70840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4469 n_71820_70840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4470 n_67260_76440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4471 n_68780_76440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4472 n_65740_79240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4473 n_64600_79240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4474 n_64600_76440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4475 n_87400_62440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4476 n_87020_59640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4477 n_88160_59640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4478 n_85880_62440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4479 n_83220_65240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4480 n_84740_62440 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4481 n_83220_68040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4482 n_84740_68040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4483 n_83600_70840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4484 n_85500_70840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4485 n_85880_68040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4486 n_85880_73640 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4487 n_81700_79240 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4488 n_85500_82040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4489 n_68780_82040 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4490 n_44460_56840 0 PWL(34000ps 0uA 34030ps 0uA 34031ps 30uA 34059ps 30uA 34060ps 0uA)
I4491 n_87020_87640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4492 n_93100_87640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4493 n_93480_56840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4494 n_90440_62440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4495 n_93100_84840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4496 n_83600_87640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4497 n_65740_40040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4498 n_56240_48440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4499 n_61940_48440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4500 n_93480_48440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4501 n_93480_54040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4502 n_63840_40040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4503 n_87020_40040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4504 n_52440_40040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4505 n_40660_42840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4506 n_42940_42840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4507 n_56620_40040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4508 n_67260_40040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4509 n_90440_40040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4510 n_93480_45640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4511 n_80560_40040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4512 n_46360_40040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4513 n_40280_40040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4514 n_72200_40040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4515 n_55100_40040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4516 n_40660_45640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4517 n_50160_59640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4518 n_43320_62440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4519 n_44460_62440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4520 n_51300_59640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4521 n_45220_48440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4522 n_54720_42840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4523 n_71820_42840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4524 n_41420_40040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4525 n_49400_40040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4526 n_80180_42840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4527 n_88920_45640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4528 n_83600_42840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4529 n_66880_45640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4530 n_57760_40040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4531 n_44840_45640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4532 n_43700_42840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4533 n_51680_42840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4534 n_87020_45640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4535 n_63460_42840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4536 n_92340_51240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4537 n_90440_48440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4538 n_60040_48440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4539 n_55100_54040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4540 n_63080_51240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4541 n_80180_87640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4542 n_90820_84840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4543 n_90820_59640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4544 n_88920_56840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4545 n_90060_87640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4546 n_85120_84840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4547 n_68780_79240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4548 n_83220_54040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4549 n_91200_54040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4550 n_92340_56840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4551 n_90820_65240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4552 n_88920_70840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4553 n_87400_65240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4554 n_92720_82040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4555 n_92340_76440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4556 n_82080_84840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4557 n_88920_87640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4558 n_83600_51240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4559 n_80560_51240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4560 n_84740_54040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4561 n_90820_56840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4562 n_77520_54040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4563 n_87400_79240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4564 n_89300_59640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4565 n_89300_73640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4566 n_92340_73640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4567 n_88920_76440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4568 n_90060_79240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4569 n_90820_82040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4570 n_77900_87640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4571 n_81700_82040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4572 n_79040_87640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4573 n_79040_54040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4574 n_80560_54040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4575 n_82080_54040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4576 n_80560_56840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4577 n_82080_56840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4578 n_78660_56840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4579 n_83600_56840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4580 n_76760_65240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4581 n_80940_62440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4582 n_76380_68040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4583 n_76000_70840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4584 n_79040_68040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4585 n_78280_70840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4586 n_75240_73640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4587 n_73720_70840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4588 n_73720_79240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4589 n_73720_73640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4590 n_70300_79240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4591 n_71820_79240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4592 n_88920_79240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4593 n_65360_87640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4594 n_72200_84840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4595 n_85500_56840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4596 n_82080_59640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4597 n_84740_65240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4598 n_83600_59640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4599 n_82080_68040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4600 n_80560_68040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4601 n_77140_70840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4602 n_79040_70840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4603 n_78660_76440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4604 n_78660_79240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4605 n_78280_82040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4606 n_76760_84840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4607 n_76380_87640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4608 n_74860_84840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4609 n_74860_82040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4610 n_76760_82040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4611 n_60800_51240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4612 n_71820_51240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4613 n_71820_54040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4614 n_53200_51240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4615 n_70300_51240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4616 n_53580_54040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4617 n_56620_51240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4618 n_68780_51240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4619 n_61940_51240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4620 n_41800_56840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4621 n_52060_51240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4622 n_70300_54040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4623 n_61560_54040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4624 n_87400_51240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4625 n_90820_51240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4626 n_65360_42840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4627 n_90440_45640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4628 n_50540_42840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4629 n_45220_42840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4630 n_46740_45640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4631 n_61560_40040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4632 n_68020_48440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4633 n_85500_42840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4634 n_88920_42840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4635 n_82080_42840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4636 n_51300_40040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4637 n_43320_40040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4638 n_73720_45640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4639 n_53200_42840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4640 n_44080_48440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4641 n_58900_48440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4642 n_48260_65240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4643 n_50920_68040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4644 n_72200_56840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4645 n_53580_59640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4646 n_53580_62440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4647 n_55100_65240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4648 n_49400_65240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4649 n_56620_65240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4650 n_61560_65240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4651 n_60420_65240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4652 n_73720_62440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4653 n_76380_62440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4654 n_76380_59640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4655 n_63080_82040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4656 n_75240_59640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4657 n_77520_62440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4658 n_73340_59640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4659 n_55100_56840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4660 n_69160_62440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4661 n_70300_73640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4662 n_56620_73640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4663 n_66880_73640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4664 n_63460_70840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4665 n_74100_68040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4666 n_65360_68040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4667 n_68780_68040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4668 n_75240_68040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4669 n_72960_68040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4670 n_63080_73640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4671 n_76760_73640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4672 n_67260_70840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4673 n_70300_48440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4674 n_41800_70840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4675 n_40660_79240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4676 n_40280_82040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4677 n_44080_84840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4678 n_40280_87640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4679 n_50920_82040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4680 n_53580_82040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4681 n_47500_56840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4682 n_44080_59640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4683 n_42940_82040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4684 n_45220_82040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4685 n_41420_87640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4686 n_46740_87640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4687 n_46740_84840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4688 n_61940_84840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4689 n_63080_84840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4690 n_49400_84840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4691 n_58140_87640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4692 n_59660_84840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4693 n_55100_82040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4694 n_46740_51240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4695 n_63080_54040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4696 n_68780_56840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4697 n_45220_87640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4698 n_59280_87640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4699 n_74860_87640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4700 n_67260_82040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4701 n_65740_82040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4702 n_53580_87640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4703 n_64600_84840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4704 n_57000_87640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4705 n_63460_59640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4706 n_63460_56840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4707 n_68780_59640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4708 n_67260_56840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4709 n_70300_59640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4710 n_70300_62440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4711 n_70300_56840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4712 n_70300_65240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4713 n_71820_65240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4714 n_71820_68040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4715 n_70300_70840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4716 n_71820_70840 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4717 n_67260_76440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4718 n_65740_79240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4719 n_64600_79240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4720 n_64600_76440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4721 n_58520_82040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4722 n_56240_82040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4723 n_84740_62440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4724 n_84740_73640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4725 n_85880_68040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4726 n_83600_76440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4727 n_85500_76440 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4728 n_85500_79240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4729 n_83600_79240 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4730 n_68780_82040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4731 n_71060_82040 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4732 n_60040_59640 0 PWL(36000ps 0uA 36030ps 0uA 36031ps 30uA 36059ps 30uA 36060ps 0uA)
I4733 n_93480_62440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4734 n_93480_79240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4735 n_91960_87640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4736 n_93480_56840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4737 n_93480_68040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4738 n_93480_73640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4739 n_93480_76440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4740 n_83600_87640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4741 n_65740_40040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4742 n_54720_48440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4743 n_65740_45640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4744 n_40280_54040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4745 n_79040_42840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4746 n_92340_48440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4747 n_41800_42840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4748 n_63840_40040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4749 n_91580_40040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4750 n_88160_40040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4751 n_52440_40040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4752 n_56620_40040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4753 n_93480_45640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4754 n_80560_40040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4755 n_40280_48440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4756 n_60040_45640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4757 n_82080_48440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4758 n_77140_40040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4759 n_43320_62440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4760 n_44460_62440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4761 n_74860_40040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4762 n_80180_45640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4763 n_56620_45640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4764 n_41420_48440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4765 n_80180_42840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4766 n_88920_45640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4767 n_57760_40040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4768 n_51680_42840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4769 n_83600_40040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4770 n_92720_40040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4771 n_63460_42840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4772 n_48260_45640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4773 n_85120_48440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4774 n_78280_48440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4775 n_47880_54040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4776 n_64600_51240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4777 n_54720_51240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4778 n_63080_51240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4779 n_80180_87640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4780 n_90440_76440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4781 n_90440_73640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4782 n_92340_65240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4783 n_88920_56840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4784 n_87400_84840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4785 n_91580_79240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4786 n_91580_62440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4787 n_68780_79240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4788 n_83220_54040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4789 n_91200_54040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4790 n_92340_56840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4791 n_88920_70840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4792 n_87400_65240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4793 n_92720_82040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4794 n_88920_82040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4795 n_88920_87640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4796 n_85880_87640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4797 n_83600_51240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4798 n_80560_51240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4799 n_84740_54040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4800 n_90820_56840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4801 n_77520_54040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4802 n_87400_79240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4803 n_88920_65240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4804 n_92340_73640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4805 n_90060_79240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4806 n_89300_84840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4807 n_90820_82040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4808 n_77900_87640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4809 n_81700_82040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4810 n_79040_87640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4811 n_79040_54040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4812 n_80560_54040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4813 n_82080_54040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4814 n_80560_56840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4815 n_82080_56840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4816 n_78660_56840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4817 n_83600_56840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4818 n_76760_65240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4819 n_80940_62440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4820 n_76760_56840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4821 n_78660_65240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4822 n_80560_65240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4823 n_77900_68040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4824 n_79040_68040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4825 n_78280_70840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4826 n_75240_76440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4827 n_70300_79240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4828 n_67260_84840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4829 n_65740_84840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4830 n_62320_82040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4831 n_68780_87640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4832 n_68780_84840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4833 n_85500_56840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4834 n_85500_59640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4835 n_84740_65240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4836 n_83600_59640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4837 n_82080_65240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4838 n_82080_68040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4839 n_82080_70840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4840 n_81700_73640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4841 n_78660_73640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4842 n_78660_76440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4843 n_78660_79240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4844 n_72200_76440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4845 n_78280_82040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4846 n_80560_79240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4847 n_76760_84840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4848 n_76380_87640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4849 n_74860_84840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4850 n_60800_51240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4851 n_71820_51240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4852 n_71820_54040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4853 n_53200_51240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4854 n_53580_54040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4855 n_68020_54040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4856 n_56620_51240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4857 n_49780_54040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4858 n_41800_56840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4859 n_52060_51240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4860 n_70300_54040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4861 n_61560_54040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4862 n_79040_51240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4863 n_83600_48440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4864 n_49400_48440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4865 n_65360_42840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4866 n_92720_42840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4867 n_85500_40040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4868 n_50540_42840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4869 n_61560_40040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4870 n_88920_42840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4871 n_82080_42840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4872 n_42940_48440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4873 n_53200_45640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4874 n_82080_45640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4875 n_73340_40040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4876 n_57000_54040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4877 n_72200_56840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4878 n_76380_62440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4879 n_75240_62440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4880 n_63080_82040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4881 n_75240_59640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4882 n_73340_59640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4883 n_75240_68040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4884 n_75240_65240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4885 n_72960_68040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4886 n_68020_62440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4887 n_68780_70840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4888 n_71820_73640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4889 n_76760_73640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4890 n_63080_79240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4891 n_61560_79240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4892 n_52060_82040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4893 n_58140_51240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4894 n_70300_48440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4895 n_41800_70840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4896 n_40660_79240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4897 n_40280_82040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4898 n_40280_87640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4899 n_57380_76440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4900 n_63080_76440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4901 n_80560_76440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4902 n_49400_82040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4903 n_54720_84840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4904 n_52820_79240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4905 n_44080_59640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4906 n_42940_82040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4907 n_45220_82040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4908 n_40280_84840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4909 n_41420_87640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4910 n_46740_87640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4911 n_63080_84840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4912 n_42940_54040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4913 n_63080_54040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4914 n_68780_56840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4915 n_67260_82040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4916 n_65740_82040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4917 n_58520_84840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4918 n_64600_84840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4919 n_73340_87640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4920 n_56240_76440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4921 n_63460_59640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4922 n_63460_56840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4923 n_68780_59640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4924 n_70300_59640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4925 n_70300_56840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4926 n_70300_65240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4927 n_71820_65240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4928 n_71820_68040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4929 n_70300_70840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4930 n_71820_70840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4931 n_67260_76440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4932 n_65740_79240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4933 n_53960_79240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4934 n_55100_79240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4935 n_58520_82040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4936 n_59660_82040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4937 n_83220_65240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4938 n_84740_62440 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4939 n_85880_68040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4940 n_83600_82040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4941 n_83600_79240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4942 n_69920_82040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4943 n_68780_82040 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4944 n_43320_65240 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4945 n_44460_56840 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4946 n_60040_59640 0 PWL(38000ps 0uA 38030ps 0uA 38031ps 30uA 38059ps 30uA 38060ps 0uA)
I4947 n_90820_68040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4948 n_91200_70840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4949 n_87020_87640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4950 n_93480_56840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4951 n_90440_62440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4952 n_93480_76440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4953 n_93100_84840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4954 n_84740_87640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4955 n_65740_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4956 n_54720_48440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4957 n_61940_48440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4958 n_40280_54040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4959 n_40660_56840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4960 n_63840_45640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4961 n_79040_42840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4962 n_92340_48440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4963 n_41800_42840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4964 n_50920_48440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4965 n_63840_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4966 n_70300_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4967 n_87020_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4968 n_40660_42840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4969 n_56620_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4970 n_67260_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4971 n_90440_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4972 n_93480_45640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4973 n_46360_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4974 n_40280_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4975 n_72200_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4976 n_79040_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4977 n_82080_48440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4978 n_77140_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4979 n_55100_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4980 n_50160_59640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4981 n_45600_68040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4982 n_40660_65240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4983 n_41800_68040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4984 n_47500_68040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4985 n_51300_59640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4986 n_54720_42840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4987 n_74860_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4988 n_80180_45640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4989 n_76760_42840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4990 n_71820_42840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4991 n_41420_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4992 n_49400_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4993 n_88920_45640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4994 n_83600_42840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4995 n_66880_45640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4996 n_57760_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4997 n_43700_42840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4998 n_87020_45640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I4999 n_68400_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5000 n_63460_42840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5001 n_51680_48440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5002 n_48260_45640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5003 n_85120_48440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5004 n_78280_48440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5005 n_64980_48440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5006 n_41420_54040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5007 n_47880_54040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5008 n_60040_48440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5009 n_54720_51240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5010 n_63080_51240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5011 n_81700_87640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5012 n_90820_84840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5013 n_90440_76440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5014 n_90820_59640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5015 n_88920_56840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5016 n_85120_84840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5017 n_87400_73640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5018 n_88540_68040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5019 n_68780_79240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5020 n_87400_65240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5021 n_87400_76440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5022 n_82080_84840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5023 n_87400_56840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5024 n_89300_59640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5025 n_88920_76440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5026 n_89300_84840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5027 n_81700_82040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5028 n_80180_59640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5029 n_82080_56840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5030 n_78660_56840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5031 n_76380_54040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5032 n_80940_62440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5033 n_76760_56840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5034 n_80560_65240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5035 n_75240_76440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5036 n_67260_84840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5037 n_71820_79240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5038 n_88920_79240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5039 n_65740_84840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5040 n_62320_82040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5041 n_70300_87640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5042 n_85500_56840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5043 n_86260_54040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5044 n_85500_59640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5045 n_84740_65240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5046 n_83600_59640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5047 n_85880_65240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5048 n_87400_68040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5049 n_81700_73640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5050 n_80560_70840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5051 n_80560_73640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5052 n_81700_76440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5053 n_72200_76440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5054 n_76760_79240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5055 n_74860_82040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5056 n_76760_82040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5057 n_67260_51240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5058 n_70300_51240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5059 n_61940_51240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5060 n_49780_54040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5061 n_52060_51240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5062 n_66120_51240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5063 n_79040_51240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5064 n_83600_48440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5065 n_49400_48440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5066 n_53200_48440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5067 n_65360_42840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5068 n_70300_42840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5069 n_90440_45640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5070 n_45220_42840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5071 n_61560_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5072 n_68020_48440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5073 n_85500_42840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5074 n_88920_42840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5075 n_51300_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5076 n_43320_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5077 n_73720_45640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5078 n_76760_45640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5079 n_82080_45640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5080 n_73340_40040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5081 n_53200_42840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5082 n_52060_54040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5083 n_48260_65240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5084 n_50920_68040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5085 n_53580_59640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5086 n_53580_62440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5087 n_55100_65240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5088 n_49400_65240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5089 n_56620_65240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5090 n_61560_65240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5091 n_60420_65240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5092 n_73720_62440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5093 n_75240_62440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5094 n_63080_82040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5095 n_75240_59640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5096 n_77520_62440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5097 n_73340_59640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5098 n_55100_56840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5099 n_69160_62440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5100 n_70300_73640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5101 n_56620_73640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5102 n_58140_79240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5103 n_63460_70840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5104 n_74100_68040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5105 n_65360_70840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5106 n_68780_68040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5107 n_75240_65240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5108 n_68020_62440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5109 n_55480_48440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5110 n_68780_70840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5111 n_47500_79240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5112 n_48640_79240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5113 n_60040_76440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5114 n_63080_73640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5115 n_71820_73640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5116 n_60040_79240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5117 n_61560_79240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5118 n_65740_76440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5119 n_46360_68040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5120 n_44840_70840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5121 n_44840_76440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5122 n_41800_70840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5123 n_40660_79240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5124 n_43700_79240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5125 n_44080_84840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5126 n_57380_76440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5127 n_63080_76440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5128 n_67260_79240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5129 n_53580_82040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5130 n_50160_84840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5131 n_70300_76440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5132 n_40280_84840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5133 n_49400_84840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5134 n_49400_87640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5135 n_64220_82040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5136 n_61940_87640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5137 n_42940_54040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5138 n_46740_51240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5139 n_43320_68040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5140 n_43320_76440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5141 n_44080_82040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5142 n_65360_56840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5143 n_63080_54040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5144 n_68780_56840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5145 n_45220_87640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5146 n_51680_84840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5147 n_54340_76440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5148 n_67260_82040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5149 n_58520_84840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5150 n_64600_84840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5151 n_73340_87640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5152 n_63460_59640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5153 n_63460_56840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5154 n_60040_54040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5155 n_68780_59640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5156 n_70300_62440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5157 n_70300_70840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5158 n_70300_68040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5159 n_71820_70840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5160 n_64600_79240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5161 n_53960_79240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5162 n_64600_76440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5163 n_56240_82040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5164 n_88160_59640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5165 n_85880_62440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5166 n_84740_62440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5167 n_85500_70840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5168 n_83220_73640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5169 n_84740_73640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5170 n_85880_68040 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5171 n_83600_76440 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5172 n_81700_79240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5173 n_43320_65240 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5174 n_60040_56840 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5175 n_60040_59640 0 PWL(40000ps 0uA 40030ps 0uA 40031ps 30uA 40059ps 30uA 40060ps 0uA)
I5176 n_91200_70840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5177 n_87020_87640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5178 n_93480_56840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5179 n_90440_62440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5180 n_93480_68040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5181 n_93480_76440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5182 n_93100_84840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5183 n_84740_87640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5184 n_65740_40040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5185 n_54720_48440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5186 n_56240_48440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5187 n_61940_48440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5188 n_63840_45640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5189 n_79040_42840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5190 n_93480_48440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5191 n_92340_48440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5192 n_63840_40040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5193 n_91580_40040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5194 n_40660_42840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5195 n_56620_40040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5196 n_67260_40040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5197 n_93480_45640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5198 n_46360_40040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5199 n_40280_40040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5200 n_60040_45640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5201 n_82080_48440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5202 n_55100_40040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5203 n_40660_45640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5204 n_40660_51240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5205 n_50160_59640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5206 n_45600_68040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5207 n_47500_68040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5208 n_51300_59640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5209 n_44840_51240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5210 n_45220_48440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5211 n_54720_42840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5212 n_80180_45640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5213 n_56620_45640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5214 n_41420_40040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5215 n_49400_40040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5216 n_88920_45640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5217 n_66880_45640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5218 n_57760_40040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5219 n_43700_42840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5220 n_92720_40040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5221 n_63460_42840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5222 n_85120_48440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5223 n_90440_48440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5224 n_78280_48440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5225 n_64980_48440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5226 n_60040_48440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5227 n_55100_54040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5228 n_54720_51240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5229 n_63080_51240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5230 n_81700_87640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5231 n_90820_84840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5232 n_90440_76440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5233 n_92340_65240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5234 n_90820_59640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5235 n_88920_56840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5236 n_85120_84840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5237 n_87400_73640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5238 n_68780_79240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5239 n_83220_54040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5240 n_91200_54040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5241 n_87400_76440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5242 n_87780_87640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5243 n_88920_82040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5244 n_82080_84840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5245 n_88920_87640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5246 n_85880_87640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5247 n_83600_51240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5248 n_80560_51240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5249 n_85500_51240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5250 n_87400_56840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5251 n_89300_59640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5252 n_88920_65240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5253 n_88920_76440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5254 n_89300_84840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5255 n_81700_82040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5256 n_80560_54040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5257 n_77900_51240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5258 n_82080_54040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5259 n_80560_56840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5260 n_80180_59640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5261 n_76380_54040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5262 n_76760_65240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5263 n_80940_62440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5264 n_76760_56840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5265 n_78660_65240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5266 n_77900_68040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5267 n_76000_70840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5268 n_78280_70840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5269 n_75240_73640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5270 n_73720_79240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5271 n_73720_73640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5272 n_67260_84840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5273 n_71820_79240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5274 n_67260_87640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5275 n_65740_84840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5276 n_62320_82040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5277 n_65360_87640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5278 n_70300_87640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5279 n_72200_84840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5280 n_82080_51240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5281 n_85500_56840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5282 n_86260_54040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5283 n_87400_48440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5284 n_85500_59640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5285 n_84740_65240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5286 n_83600_59640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5287 n_85880_65240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5288 n_77140_70840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5289 n_81700_73640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5290 n_80560_70840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5291 n_80560_73640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5292 n_81700_76440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5293 n_72200_76440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5294 n_76760_79240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5295 n_67260_51240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5296 n_71820_51240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5297 n_70300_51240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5298 n_68020_54040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5299 n_61940_51240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5300 n_75240_54040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5301 n_66120_51240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5302 n_76380_51240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5303 n_79040_51240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5304 n_87400_51240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5305 n_83600_48440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5306 n_65360_42840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5307 n_92720_42840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5308 n_45220_42840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5309 n_61560_40040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5310 n_68020_48440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5311 n_88920_42840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5312 n_51300_40040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5313 n_43320_40040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5314 n_53200_45640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5315 n_82080_45640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5316 n_53200_42840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5317 n_44080_48440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5318 n_43320_51240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5319 n_57000_54040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5320 n_52060_54040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5321 n_48260_65240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5322 n_50920_68040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5323 n_72200_56840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5324 n_53580_59640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5325 n_53580_62440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5326 n_55100_65240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5327 n_49400_65240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5328 n_56620_65240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5329 n_61560_62440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5330 n_58520_65240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5331 n_59660_68040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5332 n_60800_68040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5333 n_60040_73640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5334 n_63080_65240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5335 n_76380_59640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5336 n_63080_82040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5337 n_72200_62440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5338 n_73340_59640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5339 n_61940_68040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5340 n_59660_70840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5341 n_50920_73640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5342 n_49400_73640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5343 n_55860_68040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5344 n_49780_76440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5345 n_50920_79240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5346 n_61560_73640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5347 n_58520_73640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5348 n_70300_73640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5349 n_66880_73640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5350 n_65360_68040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5351 n_65360_70840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5352 n_47500_79240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5353 n_48640_79240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5354 n_60040_76440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5355 n_63080_73640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5356 n_71820_73640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5357 n_56620_79240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5358 n_52060_82040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5359 n_67260_70840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5360 n_58140_51240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5361 n_70300_48440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5362 n_46360_68040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5363 n_44840_70840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5364 n_44840_76440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5365 n_41800_70840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5366 n_40660_79240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5367 n_43700_79240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5368 n_40280_87640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5369 n_57380_76440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5370 n_63080_76440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5371 n_67260_79240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5372 n_50920_82040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5373 n_50160_84840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5374 n_65740_73640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5375 n_70300_76440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5376 n_47500_56840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5377 n_52820_79240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5378 n_40280_84840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5379 n_41420_87640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5380 n_46740_87640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5381 n_46740_84840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5382 n_52440_87640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5383 n_49400_87640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5384 n_64220_82040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5385 n_58140_87640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5386 n_55100_82040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5387 n_61940_87640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5388 n_65360_59640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5389 n_54340_76440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5390 n_54340_87640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5391 n_67260_82040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5392 n_53580_87640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5393 n_58520_84840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5394 n_64600_84840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5395 n_57000_87640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5396 n_65360_65240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5397 n_63460_62440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5398 n_70300_59640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5399 n_70300_62440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5400 n_70300_56840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5401 n_71820_59640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5402 n_70300_65240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5403 n_71820_65240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5404 n_71820_68040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5405 n_70300_68040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5406 n_67260_76440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5407 n_68780_76440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5408 n_65740_79240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5409 n_64600_79240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5410 n_64600_76440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5411 n_87400_62440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5412 n_88920_62440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5413 n_83220_62440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5414 n_83220_68040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5415 n_84740_68040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5416 n_83600_70840 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5417 n_83220_73640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5418 n_85880_73640 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5419 n_85500_76440 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5420 n_85500_79240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5421 n_83600_82040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5422 n_69920_82040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5423 n_71060_82040 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5424 n_43320_65240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5425 n_75240_51240 0 PWL(42000ps 0uA 42030ps 0uA 42031ps 30uA 42059ps 30uA 42060ps 0uA)
I5426 n_93480_62440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5427 n_91960_87640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5428 n_93100_87640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5429 n_93480_56840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5430 n_93480_73640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5431 n_83600_87640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5432 n_84740_87640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5433 n_54720_48440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5434 n_79040_42840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5435 n_70300_40040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5436 n_91580_40040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5437 n_87020_40040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5438 n_88160_40040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5439 n_52440_40040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5440 n_40660_42840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5441 n_67260_40040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5442 n_93480_45640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5443 n_80560_40040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5444 n_46360_40040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5445 n_40280_48440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5446 n_60040_45640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5447 n_82080_48440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5448 n_77140_40040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5449 n_40660_45640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5450 n_50160_59640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5451 n_42180_73640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5452 n_44460_68040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5453 n_46740_65240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5454 n_52060_73640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5455 n_51300_59640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5456 n_45220_48440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5457 n_74860_40040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5458 n_80180_45640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5459 n_56620_45640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5460 n_41420_48440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5461 n_49400_40040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5462 n_80180_42840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5463 n_88920_45640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5464 n_66880_45640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5465 n_43700_42840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5466 n_51680_42840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5467 n_83600_40040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5468 n_87020_45640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5469 n_92720_40040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5470 n_68400_40040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5471 n_78280_48440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5472 n_54720_51240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5473 n_81700_87640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5474 n_80180_87640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5475 n_90440_73640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5476 n_88920_56840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5477 n_90060_87640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5478 n_87400_84840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5479 n_91580_62440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5480 n_92340_56840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5481 n_87780_87640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5482 n_88920_87640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5483 n_84740_54040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5484 n_90820_56840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5485 n_77520_54040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5486 n_87400_79240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5487 n_92340_73640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5488 n_89300_84840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5489 n_90820_82040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5490 n_77900_87640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5491 n_81700_82040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5492 n_79040_54040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5493 n_77900_51240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5494 n_83600_56840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5495 n_76760_65240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5496 n_80940_62440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5497 n_76760_56840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5498 n_78660_65240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5499 n_77900_68040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5500 n_76000_70840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5501 n_75240_73640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5502 n_73720_79240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5503 n_73720_73640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5504 n_70300_79240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5505 n_67260_84840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5506 n_67260_87640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5507 n_65740_84840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5508 n_62320_82040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5509 n_65360_87640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5510 n_68780_87640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5511 n_68780_84840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5512 n_70300_87640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5513 n_72200_84840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5514 n_85500_56840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5515 n_85500_59640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5516 n_87400_68040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5517 n_80560_68040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5518 n_80560_70840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5519 n_80560_73640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5520 n_76760_76440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5521 n_80560_79240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5522 n_71820_51240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5523 n_70300_51240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5524 n_75240_54040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5525 n_76380_51240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5526 n_79040_51240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5527 n_70300_42840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5528 n_92720_42840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5529 n_90440_45640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5530 n_85500_40040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5531 n_50540_42840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5532 n_45220_42840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5533 n_68020_48440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5534 n_88920_42840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5535 n_82080_42840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5536 n_51300_40040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5537 n_42940_48440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5538 n_53200_45640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5539 n_82080_45640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5540 n_73340_40040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5541 n_44080_48440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5542 n_58900_48440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5543 n_58520_59640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5544 n_52060_54040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5545 n_48260_65240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5546 n_50920_68040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5547 n_51680_62440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5548 n_49400_65240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5549 n_56620_65240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5550 n_58520_65240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5551 n_60420_65240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5552 n_73720_62440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5553 n_75240_62440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5554 n_76380_59640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5555 n_58140_62440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5556 n_53580_73640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5557 n_46360_76440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5558 n_48260_73640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5559 n_61560_73640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5560 n_66880_73640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5561 n_56620_70840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5562 n_68780_70840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5563 n_46740_62440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5564 n_46740_70840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5565 n_48260_76440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5566 n_47500_79240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5567 n_45600_84840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5568 n_48640_79240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5569 n_58520_70840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5570 n_60040_76440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5571 n_60420_70840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5572 n_63080_73640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5573 n_56620_79240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5574 n_65740_76440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5575 n_67260_70840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5576 n_58140_51240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5577 n_56620_62440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5578 n_70300_48440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5579 n_41800_70840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5580 n_40660_79240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5581 n_40280_82040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5582 n_44080_84840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5583 n_57380_76440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5584 n_80560_76440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5585 n_49400_82040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5586 n_54720_84840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5587 n_65740_73640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5588 n_47500_56840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5589 n_40280_84840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5590 n_41420_87640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5591 n_46740_87640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5592 n_43320_87640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5593 n_61940_84840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5594 n_42940_54040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5595 n_65360_59640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5596 n_65360_56840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5597 n_68780_56840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5598 n_59280_87640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5599 n_60800_84840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5600 n_61180_82040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5601 n_54340_76440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5602 n_67260_56840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5603 n_71820_59640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5604 n_71820_70840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5605 n_68780_76440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5606 n_55100_79240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5607 n_87020_59640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5608 n_83220_62440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5609 n_83220_68040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5610 n_84740_68040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5611 n_83600_70840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5612 n_85500_70840 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5613 n_83220_73640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5614 n_84740_73640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5615 n_85880_73640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5616 n_83600_76440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5617 n_81700_79240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5618 n_85500_76440 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5619 n_85500_79240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5620 n_83600_82040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5621 n_69920_82040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5622 n_71060_82040 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5623 n_43320_65240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5624 n_60040_59640 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5625 n_75240_51240 0 PWL(44000ps 0uA 44030ps 0uA 44031ps 30uA 44059ps 30uA 44060ps 0uA)
I5626 n_92340_54040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5627 n_93480_62440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5628 n_93480_79240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5629 n_93480_73640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5630 n_93480_76440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5631 n_93100_84840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5632 n_83600_87640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5633 n_65740_40040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5634 n_54720_48440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5635 n_61940_48440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5636 n_63840_45640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5637 n_79040_42840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5638 n_92340_48440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5639 n_91580_40040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5640 n_87020_40040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5641 n_88160_40040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5642 n_52440_40040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5643 n_56620_40040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5644 n_67260_40040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5645 n_46360_40040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5646 n_40280_48440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5647 n_82080_48440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5648 n_77140_40040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5649 n_40660_51240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5650 n_42180_73640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5651 n_44460_68040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5652 n_46740_65240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5653 n_52060_73640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5654 n_44840_51240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5655 n_74860_40040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5656 n_80180_45640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5657 n_41420_48440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5658 n_49400_40040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5659 n_66880_45640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5660 n_57760_40040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5661 n_51680_42840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5662 n_83600_40040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5663 n_87020_45640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5664 n_92720_40040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5665 n_85120_48440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5666 n_78280_48440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5667 n_64980_48440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5668 n_60040_48440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5669 n_54720_51240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5670 n_63080_51240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5671 n_80180_87640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5672 n_90820_84840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5673 n_90440_76440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5674 n_90440_73640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5675 n_91580_79240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5676 n_91580_62440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5677 n_89300_54040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5678 n_68780_79240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5679 n_88920_51240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5680 n_83220_54040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5681 n_91200_54040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5682 n_92340_56840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5683 n_92340_76440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5684 n_83600_51240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5685 n_80560_51240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5686 n_85500_51240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5687 n_84740_54040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5688 n_87400_56840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5689 n_90820_56840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5690 n_77520_54040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5691 n_87400_79240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5692 n_92340_73640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5693 n_88920_76440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5694 n_90820_82040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5695 n_77900_87640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5696 n_79040_54040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5697 n_80560_54040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5698 n_82080_54040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5699 n_80560_56840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5700 n_82080_56840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5701 n_78660_56840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5702 n_83600_56840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5703 n_76380_54040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5704 n_80940_62440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5705 n_76760_56840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5706 n_76380_68040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5707 n_78280_70840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5708 n_70300_79240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5709 n_71820_79240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5710 n_71820_87640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5711 n_82080_51240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5712 n_85500_56840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5713 n_85500_59640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5714 n_87400_68040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5715 n_80560_68040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5716 n_80560_70840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5717 n_80560_73640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5718 n_76760_76440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5719 n_72200_76440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5720 n_74860_84840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5721 n_74860_82040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5722 n_76760_82040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5723 n_67260_51240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5724 n_70300_51240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5725 n_61940_51240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5726 n_66120_51240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5727 n_79040_51240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5728 n_83600_48440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5729 n_92720_42840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5730 n_90440_45640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5731 n_85500_40040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5732 n_50540_42840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5733 n_61560_40040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5734 n_68020_48440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5735 n_51300_40040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5736 n_42940_48440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5737 n_82080_45640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5738 n_73340_40040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5739 n_43320_51240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5740 n_58520_59640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5741 n_48260_65240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5742 n_49780_62440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5743 n_59660_62440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5744 n_44840_73640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5745 n_50920_68040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5746 n_51680_62440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5747 n_53580_59640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5748 n_53580_62440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5749 n_52060_65240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5750 n_56620_65240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5751 n_58520_65240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5752 n_60420_65240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5753 n_73720_62440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5754 n_75240_62440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5755 n_76380_59640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5756 n_63080_82040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5757 n_72200_62440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5758 n_73340_59640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5759 n_55100_56840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5760 n_58140_62440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5761 n_69160_62440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5762 n_53580_73640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5763 n_50920_73640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5764 n_46740_73640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5765 n_40660_76440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5766 n_40660_70840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5767 n_65360_68040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5768 n_65360_70840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5769 n_56620_70840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5770 n_46740_62440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5771 n_46740_70840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5772 n_45600_84840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5773 n_71820_73640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5774 n_76760_73640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5775 n_56620_79240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5776 n_60040_79240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5777 n_63080_79240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5778 n_65740_76440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5779 n_56620_62440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5780 n_41800_70840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5781 n_43700_79240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5782 n_57380_76440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5783 n_63080_76440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5784 n_50920_82040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5785 n_53580_82040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5786 n_70300_76440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5787 n_47500_56840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5788 n_52820_79240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5789 n_41420_87640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5790 n_46740_87640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5791 n_43320_87640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5792 n_46740_84840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5793 n_61940_84840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5794 n_63080_84840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5795 n_49400_84840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5796 n_52440_87640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5797 n_58140_87640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5798 n_55100_82040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5799 n_65360_62440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5800 n_66880_62440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5801 n_65360_56840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5802 n_68780_56840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5803 n_45220_87640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5804 n_59280_87640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5805 n_51680_84840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5806 n_60800_84840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5807 n_61180_82040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5808 n_54340_76440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5809 n_54340_87640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5810 n_67260_82040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5811 n_65740_82040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5812 n_53580_87640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5813 n_58520_84840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5814 n_64600_84840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5815 n_57000_87640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5816 n_67260_65240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5817 n_63460_62440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5818 n_67260_56840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5819 n_66880_59640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5820 n_71820_59640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5821 n_68400_65240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5822 n_71820_65240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5823 n_71820_68040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5824 n_70300_70840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5825 n_67260_76440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5826 n_65740_79240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5827 n_64600_79240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5828 n_64600_76440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5829 n_55100_79240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5830 n_83220_62440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5831 n_83220_68040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5832 n_83600_70840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5833 n_85500_70840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5834 n_83220_73640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5835 n_84740_73640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5836 n_83600_76440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5837 n_85500_76440 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5838 n_85500_79240 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5839 n_83600_82040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5840 n_69920_82040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5841 n_68780_82040 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5842 n_44460_56840 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5843 n_60040_59640 0 PWL(46000ps 0uA 46030ps 0uA 46031ps 30uA 46059ps 30uA 46060ps 0uA)
I5844 n_92340_54040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5845 n_93480_62440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5846 n_91200_70840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5847 n_91960_87640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5848 n_93100_87640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5849 n_93480_56840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5850 n_90440_62440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5851 n_93480_73640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5852 n_83600_87640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5853 n_65740_40040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5854 n_54720_48440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5855 n_65740_45640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5856 n_44080_54040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5857 n_63840_45640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5858 n_79040_42840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5859 n_93480_54040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5860 n_48640_40040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5861 n_63840_40040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5862 n_70300_40040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5863 n_91580_40040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5864 n_87020_40040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5865 n_52440_40040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5866 n_93480_45640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5867 n_80560_40040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5868 n_46360_40040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5869 n_40280_40040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5870 n_40280_48440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5871 n_60040_45640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5872 n_79040_40040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5873 n_82080_48440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5874 n_77140_40040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5875 n_55100_40040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5876 n_43320_59640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5877 n_50160_59640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5878 n_51300_59640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5879 n_46740_59640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5880 n_54720_42840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5881 n_74860_40040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5882 n_80180_45640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5883 n_76760_42840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5884 n_56620_45640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5885 n_41420_48440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5886 n_41420_40040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5887 n_49400_40040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5888 n_80180_42840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5889 n_88920_45640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5890 n_51680_42840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5891 n_87020_45640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5892 n_92720_40040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5893 n_68400_40040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5894 n_63460_42840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5895 n_47880_42840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5896 n_92340_51240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5897 n_78280_48440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5898 n_64980_48440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5899 n_49020_51240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5900 n_64600_51240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5901 n_54720_51240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5902 n_63080_51240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5903 n_80180_87640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5904 n_90440_73640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5905 n_90820_59640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5906 n_88920_56840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5907 n_90060_87640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5908 n_87400_84840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5909 n_87400_73640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5910 n_91580_62440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5911 n_89300_54040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5912 n_68780_79240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5913 n_88920_51240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5914 n_90820_65240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5915 n_87400_76440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5916 n_88920_82040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5917 n_85880_87640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5918 n_87400_56840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5919 n_89300_59640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5920 n_89300_73640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5921 n_80560_84840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5922 n_76380_54040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5923 n_76760_56840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5924 n_78660_65240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5925 n_77900_68040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5926 n_76000_70840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5927 n_75240_73640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5928 n_73720_70840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5929 n_73720_79240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5930 n_73720_73640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5931 n_65360_87640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5932 n_71820_87640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5933 n_70300_87640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5934 n_70300_84840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5935 n_73720_82040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5936 n_72200_84840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5937 n_87400_48440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5938 n_82080_59640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5939 n_85500_59640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5940 n_82080_65240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5941 n_80560_73640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5942 n_78280_82040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5943 n_76760_79240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5944 n_80560_79240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5945 n_80180_82040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5946 n_74860_84840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5947 n_67260_51240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5948 n_70300_51240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5949 n_68780_51240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5950 n_50920_51240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5951 n_66120_51240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5952 n_79040_51240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5953 n_90820_51240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5954 n_51680_45640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5955 n_65360_42840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5956 n_70300_42840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5957 n_92720_42840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5958 n_90440_45640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5959 n_50540_42840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5960 n_88920_42840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5961 n_82080_42840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5962 n_51300_40040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5963 n_43320_40040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5964 n_42940_48440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5965 n_53200_45640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5966 n_76760_45640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5967 n_82080_45640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5968 n_73340_40040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5969 n_53200_42840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5970 n_58900_48440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5971 n_57000_54040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5972 n_49780_56840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5973 n_48260_62440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5974 n_48260_65240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5975 n_50920_68040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5976 n_53580_59640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5977 n_53580_62440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5978 n_52060_65240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5979 n_49400_65240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5980 n_56620_65240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5981 n_58520_65240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5982 n_60420_65240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5983 n_73720_62440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5984 n_75240_62440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5985 n_76380_59640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5986 n_63080_82040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5987 n_77520_62440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5988 n_72200_62440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5989 n_73340_59640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5990 n_69160_62440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5991 n_61560_73640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5992 n_58520_73640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5993 n_70300_73640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5994 n_66880_73640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5995 n_65360_68040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5996 n_65360_70840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5997 n_68780_70840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5998 n_63080_73640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I5999 n_76760_73640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6000 n_67260_70840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6001 n_70300_48440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6002 n_65740_73640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6003 n_70300_76440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6004 n_61940_84840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6005 n_63080_84840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6006 n_52440_87640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6007 n_49400_87640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6008 n_64220_82040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6009 n_58140_87640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6010 n_66880_62440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6011 n_65360_54040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6012 n_63080_54040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6013 n_54340_87640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6014 n_65740_82040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6015 n_53580_87640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6016 n_58520_84840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6017 n_64600_84840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6018 n_57000_87640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6019 n_67260_65240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6020 n_63460_62440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6021 n_60040_54040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6022 n_66880_59640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6023 n_71820_59640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6024 n_68400_65240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6025 n_71820_65240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6026 n_71820_68040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6027 n_70300_70840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6028 n_67260_76440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6029 n_65740_79240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6030 n_64600_79240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6031 n_64600_76440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6032 n_59660_82040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6033 n_87400_62440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6034 n_88920_62440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6035 n_87020_59640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6036 n_88160_59640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6037 n_85880_62440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6038 n_83220_65240 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6039 n_84740_62440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6040 n_83220_62440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6041 n_83220_68040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6042 n_83600_70840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6043 n_85500_70840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6044 n_83220_73640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6045 n_84740_73640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6046 n_83600_76440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6047 n_85500_76440 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6048 n_87400_82040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6049 n_71060_82040 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6050 n_60040_56840 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6051 n_60040_59640 0 PWL(48000ps 0uA 48030ps 0uA 48031ps 30uA 48059ps 30uA 48060ps 0uA)
I6052 n_92340_54040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6053 n_93480_62440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6054 n_91960_87640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6055 n_87020_87640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6056 n_93480_56840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6057 n_93480_68040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6058 n_93480_76440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6059 n_83600_87640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6060 n_65740_45640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6061 n_61940_48440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6062 n_40660_56840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6063 n_63840_45640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6064 n_79040_42840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6065 n_50920_48440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6066 n_63840_40040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6067 n_87020_40040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6068 n_88160_40040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6069 n_42940_42840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6070 n_56620_40040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6071 n_67260_40040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6072 n_90440_40040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6073 n_93480_45640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6074 n_80560_40040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6075 n_46360_40040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6076 n_40280_40040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6077 n_40280_48440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6078 n_72200_40040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6079 n_77140_40040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6080 n_40660_45640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6081 n_40660_51240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6082 n_43320_62440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6083 n_40660_65240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6084 n_41800_68040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6085 n_44460_62440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6086 n_44840_51240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6087 n_45220_48440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6088 n_74860_40040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6089 n_71820_42840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6090 n_41420_48440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6091 n_41420_40040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6092 n_49400_40040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6093 n_80180_42840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6094 n_88920_45640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6095 n_83600_42840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6096 n_66880_45640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6097 n_57760_40040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6098 n_44840_45640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6099 n_83600_40040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6100 n_87020_45640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6101 n_63460_42840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6102 n_51680_48440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6103 n_78280_48440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6104 n_64980_48440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6105 n_41420_54040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6106 n_60040_48440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6107 n_64600_51240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6108 n_80180_87640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6109 n_90440_76440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6110 n_92340_65240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6111 n_88920_56840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6112 n_85120_84840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6113 n_87400_84840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6114 n_91580_62440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6115 n_89300_54040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6116 n_87780_54040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6117 n_83220_54040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6118 n_91200_54040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6119 n_90820_65240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6120 n_87400_70840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6121 n_87400_76440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6122 n_92720_82040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6123 n_92340_76440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6124 n_88920_82040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6125 n_83600_84840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6126 n_88920_87640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6127 n_85880_87640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6128 n_83600_51240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6129 n_80560_51240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6130 n_84740_54040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6131 n_90820_56840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6132 n_77520_54040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6133 n_87400_79240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6134 n_89300_59640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6135 n_92720_59640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6136 n_91960_68040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6137 n_89300_73640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6138 n_92340_73640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6139 n_88920_76440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6140 n_80560_84840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6141 n_79040_54040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6142 n_80560_54040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6143 n_82080_54040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6144 n_76380_54040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6145 n_76760_56840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6146 n_78660_65240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6147 n_80560_65240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6148 n_67260_84840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6149 n_67260_87640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6150 n_68780_87640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6151 n_68780_84840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6152 n_85500_56840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6153 n_87400_48440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6154 n_82080_59640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6155 n_84740_65240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6156 n_82080_65240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6157 n_82080_68040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6158 n_82080_70840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6159 n_81700_73640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6160 n_78660_73640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6161 n_78660_76440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6162 n_78660_79240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6163 n_76760_79240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6164 n_80560_79240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6165 n_80180_82040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6166 n_76760_84840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6167 n_76380_87640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6168 n_74860_84840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6169 n_76760_82040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6170 n_71820_51240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6171 n_71820_54040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6172 n_53200_51240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6173 n_70300_51240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6174 n_68780_51240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6175 n_61940_51240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6176 n_47880_51240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6177 n_50920_51240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6178 n_41800_56840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6179 n_70300_54040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6180 n_61560_54040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6181 n_66120_51240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6182 n_79040_51240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6183 n_53200_48440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6184 n_65360_42840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6185 n_90440_45640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6186 n_85500_40040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6187 n_46740_45640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6188 n_61560_40040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6189 n_68020_48440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6190 n_85500_42840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6191 n_88920_42840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6192 n_82080_42840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6193 n_51300_40040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6194 n_43320_40040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6195 n_42940_48440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6196 n_73720_45640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6197 n_73340_40040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6198 n_44080_48440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6199 n_43320_51240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6200 n_61940_59640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6201 n_48260_62440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6202 n_51680_56840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6203 n_52060_54040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6204 n_49780_62440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6205 n_59660_62440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6206 n_44840_73640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6207 n_72200_56840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6208 n_49400_65240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6209 n_75240_59640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6210 n_72200_62440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6211 n_55100_56840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6212 n_50920_73640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6213 n_46740_73640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6214 n_40660_76440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6215 n_40660_70840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6216 n_46740_70840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6217 n_58140_51240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6218 n_41800_70840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6219 n_40280_82040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6220 n_40280_87640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6221 n_50920_82040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6222 n_53580_82040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6223 n_47500_56840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6224 n_52820_79240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6225 n_44080_59640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6226 n_42940_56840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6227 n_40280_84840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6228 n_41420_87640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6229 n_46740_87640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6230 n_46740_84840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6231 n_49400_84840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6232 n_55100_82040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6233 n_43320_68040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6234 n_44080_65240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6235 n_65360_62440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6236 n_65360_54040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6237 n_65360_56840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6238 n_74860_87640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6239 n_66880_59640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6240 n_71820_59640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6241 n_55100_79240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6242 n_87400_62440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6243 n_87020_59640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6244 n_88160_59640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6245 n_83220_65240 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6246 n_85500_70840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6247 n_84740_73640 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6248 n_83600_76440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6249 n_85500_76440 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6250 n_87400_82040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6251 n_85500_82040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6252 n_68780_82040 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6253 n_61560_56840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6254 n_44460_56840 0 PWL(50000ps 0uA 50030ps 0uA 50031ps 30uA 50059ps 30uA 50060ps 0uA)
I6255 n_92340_54040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6256 n_93480_79240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6257 n_91960_87640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6258 n_87020_87640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6259 n_93100_87640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6260 n_90440_62440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6261 n_93480_68040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6262 n_54720_48440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6263 n_65740_45640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6264 n_61940_48440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6265 n_40280_54040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6266 n_44080_54040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6267 n_63840_45640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6268 n_92340_48440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6269 n_41800_42840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6270 n_48640_40040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6271 n_50920_48440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6272 n_63840_40040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6273 n_91580_40040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6274 n_87020_40040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6275 n_52440_40040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6276 n_40660_42840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6277 n_67260_40040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6278 n_90440_40040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6279 n_40280_40040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6280 n_40280_48440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6281 n_60040_45640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6282 n_79040_40040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6283 n_77140_40040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6284 n_55100_40040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6285 n_40660_45640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6286 n_40660_51240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6287 n_43320_59640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6288 n_44460_68040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6289 n_43320_62440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6290 n_40660_65240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6291 n_41800_68040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6292 n_44460_62440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6293 n_46740_65240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6294 n_46740_59640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6295 n_44840_51240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6296 n_45220_48440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6297 n_54720_42840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6298 n_74860_40040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6299 n_76760_42840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6300 n_56620_45640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6301 n_41420_48440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6302 n_41420_40040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6303 n_83600_42840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6304 n_66880_45640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6305 n_43700_42840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6306 n_51680_42840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6307 n_87020_45640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6308 n_92720_40040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6309 n_63460_42840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6310 n_51680_48440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6311 n_47880_42840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6312 n_48260_45640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6313 n_85120_48440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6314 n_64980_48440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6315 n_49020_51240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6316 n_47880_54040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6317 n_60040_48440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6318 n_64600_51240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6319 n_54720_51240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6320 n_92340_65240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6321 n_90820_59640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6322 n_90060_87640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6323 n_85120_84840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6324 n_87400_84840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6325 n_91580_79240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6326 n_89300_54040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6327 n_68780_79240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6328 n_87780_54040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6329 n_92720_82040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6330 n_87780_87640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6331 n_83600_84840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6332 n_88920_87640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6333 n_92720_59640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6334 n_91960_68040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6335 n_80560_56840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6336 n_82080_56840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6337 n_78660_56840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6338 n_83600_56840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6339 n_76380_54040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6340 n_76760_65240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6341 n_76380_68040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6342 n_78660_65240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6343 n_80560_65240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6344 n_78280_70840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6345 n_71820_79240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6346 n_65740_84840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6347 n_62320_82040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6348 n_70300_87640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6349 n_70300_84840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6350 n_73720_82040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6351 n_87400_48440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6352 n_80560_73640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6353 n_79040_70840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6354 n_72200_76440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6355 n_78660_84840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6356 n_76380_87640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6357 n_76760_82040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6358 n_53200_51240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6359 n_56620_51240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6360 n_59280_51240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6361 n_46360_54040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6362 n_47880_51240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6363 n_66120_51240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6364 n_83600_48440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6365 n_49400_48440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6366 n_51680_45640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6367 n_53200_48440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6368 n_65360_42840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6369 n_92720_42840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6370 n_90440_45640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6371 n_50540_42840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6372 n_45220_42840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6373 n_68020_48440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6374 n_85500_42840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6375 n_43320_40040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6376 n_42940_48440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6377 n_53200_45640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6378 n_76760_45640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6379 n_73340_40040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6380 n_53200_42840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6381 n_44080_48440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6382 n_43320_51240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6383 n_58900_48440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6384 n_61940_59640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6385 n_49780_56840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6386 n_51680_56840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6387 n_52060_54040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6388 n_48260_65240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6389 n_59660_62440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6390 n_50920_68040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6391 n_49400_65240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6392 n_56620_65240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6393 n_58520_65240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6394 n_60420_65240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6395 n_73720_62440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6396 n_63460_68040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6397 n_75240_62440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6398 n_76380_59640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6399 n_63080_82040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6400 n_75240_59640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6401 n_77520_62440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6402 n_73340_59640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6403 n_50920_73640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6404 n_49400_73640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6405 n_55860_68040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6406 n_46360_76440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6407 n_40660_76440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6408 n_48260_73640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6409 n_40660_70840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6410 n_49780_76440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6411 n_50920_79240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6412 n_58520_68040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6413 n_61560_73640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6414 n_58520_73640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6415 n_70300_73640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6416 n_66880_73640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6417 n_63460_70840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6418 n_65360_68040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6419 n_68780_68040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6420 n_72960_68040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6421 n_55480_48440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6422 n_68780_70840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6423 n_53580_65240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6424 n_53580_68040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6425 n_49400_70840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6426 n_48260_76440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6427 n_45600_84840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6428 n_48640_79240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6429 n_49400_79240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6430 n_60040_76440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6431 n_63080_73640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6432 n_76760_73640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6433 n_60040_79240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6434 n_63080_79240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6435 n_67260_70840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6436 n_58140_51240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6437 n_41800_70840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6438 n_40280_82040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6439 n_40280_87640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6440 n_67260_79240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6441 n_80560_76440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6442 n_65740_73640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6443 n_70300_76440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6444 n_47500_56840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6445 n_52820_79240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6446 n_44080_59640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6447 n_42940_56840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6448 n_40280_84840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6449 n_43320_87640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6450 n_61940_84840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6451 n_63080_84840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6452 n_49400_87640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6453 n_64220_82040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6454 n_55100_82040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6455 n_61940_87640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6456 n_42940_54040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6457 n_43320_68040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6458 n_44080_65240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6459 n_65360_62440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6460 n_66880_62440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6461 n_63080_54040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6462 n_68780_56840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6463 n_45220_87640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6464 n_59280_87640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6465 n_51680_84840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6466 n_60800_84840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6467 n_60800_87640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6468 n_54340_76440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6469 n_65740_82040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6470 n_58520_84840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6471 n_64600_84840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6472 n_57000_87640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6473 n_63460_87640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6474 n_67260_65240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6475 n_63460_62440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6476 n_60040_54040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6477 n_68780_59640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6478 n_67260_56840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6479 n_66880_59640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6480 n_70300_59640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6481 n_70300_56840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6482 n_71820_59640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6483 n_70300_65240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6484 n_71820_65240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6485 n_73720_65240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6486 n_68780_76440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6487 n_65740_79240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6488 n_53960_79240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6489 n_55100_79240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6490 n_59660_82040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6491 n_85880_62440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6492 n_84740_62440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6493 n_83220_62440 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6494 n_83220_68040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6495 n_84740_68040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6496 n_83600_70840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6497 n_83220_73640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6498 n_81700_79240 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6499 n_68780_82040 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6500 n_61560_56840 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6501 n_60040_59640 0 PWL(52000ps 0uA 52030ps 0uA 52031ps 30uA 52059ps 30uA 52060ps 0uA)
I6502 n_92340_54040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6503 n_90820_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6504 n_91200_70840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6505 n_87020_87640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6506 n_93480_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6507 n_93480_73640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6508 n_93100_84840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6509 n_84740_87640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6510 n_65740_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6511 n_56240_48440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6512 n_65740_45640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6513 n_40660_56840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6514 n_63840_45640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6515 n_93480_48440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6516 n_93480_54040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6517 n_50920_48440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6518 n_63840_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6519 n_91580_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6520 n_87020_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6521 n_88160_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6522 n_40660_42840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6523 n_56620_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6524 n_46360_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6525 n_40280_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6526 n_40280_48440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6527 n_60040_45640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6528 n_72200_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6529 n_79040_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6530 n_82080_48440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6531 n_77140_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6532 n_55100_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6533 n_40660_45640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6534 n_50160_59640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6535 n_43320_62440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6536 n_40660_65240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6537 n_41800_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6538 n_44460_62440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6539 n_51300_59640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6540 n_45220_48440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6541 n_54720_42840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6542 n_74860_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6543 n_80180_45640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6544 n_76760_42840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6545 n_71820_42840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6546 n_56620_45640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6547 n_41420_48440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6548 n_41420_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6549 n_49400_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6550 n_57760_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6551 n_43700_42840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6552 n_83600_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6553 n_87020_45640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6554 n_92720_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6555 n_63460_42840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6556 n_51680_48440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6557 n_92340_51240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6558 n_90440_48440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6559 n_64980_48440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6560 n_41420_54040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6561 n_64600_51240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6562 n_55100_54040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6563 n_63080_51240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6564 n_81700_87640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6565 n_90820_84840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6566 n_90440_73640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6567 n_92340_65240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6568 n_85120_84840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6569 n_87400_73640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6570 n_88540_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6571 n_89300_54040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6572 n_88920_51240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6573 n_83220_54040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6574 n_91200_54040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6575 n_87400_65240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6576 n_87400_70840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6577 n_87780_87640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6578 n_88920_82040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6579 n_82080_84840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6580 n_83600_51240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6581 n_80560_51240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6582 n_84740_54040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6583 n_87400_56840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6584 n_90820_56840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6585 n_77520_54040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6586 n_87400_79240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6587 n_88920_65240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6588 n_92340_73640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6589 n_89300_84840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6590 n_81700_82040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6591 n_79040_54040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6592 n_80560_54040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6593 n_82080_54040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6594 n_80560_56840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6595 n_80180_59640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6596 n_82080_56840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6597 n_78660_56840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6598 n_83600_56840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6599 n_76380_54040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6600 n_76760_65240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6601 n_78660_65240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6602 n_77900_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6603 n_76000_70840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6604 n_78280_70840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6605 n_75240_73640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6606 n_73720_70840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6607 n_73720_79240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6608 n_73720_73640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6609 n_70300_87640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6610 n_85500_56840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6611 n_87400_48440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6612 n_85500_59640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6613 n_84740_65240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6614 n_82080_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6615 n_87400_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6616 n_82080_70840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6617 n_77140_70840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6618 n_81700_73640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6619 n_78660_73640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6620 n_79040_70840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6621 n_78660_76440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6622 n_78660_79240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6623 n_78280_82040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6624 n_80560_79240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6625 n_76760_84840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6626 n_78660_84840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6627 n_74860_84840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6628 n_74860_82040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6629 n_76760_82040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6630 n_60800_51240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6631 n_53580_54040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6632 n_56620_51240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6633 n_41800_56840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6634 n_66120_51240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6635 n_87400_51240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6636 n_90820_51240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6637 n_53200_48440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6638 n_65360_42840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6639 n_92720_42840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6640 n_90440_45640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6641 n_85500_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6642 n_45220_42840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6643 n_61560_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6644 n_51300_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6645 n_43320_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6646 n_42940_48440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6647 n_53200_45640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6648 n_73720_45640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6649 n_76760_45640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6650 n_82080_45640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6651 n_73340_40040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6652 n_53200_42840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6653 n_44080_48440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6654 n_57000_54040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6655 n_48260_65240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6656 n_50920_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6657 n_72200_56840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6658 n_53580_59640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6659 n_53580_62440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6660 n_52060_65240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6661 n_49400_65240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6662 n_56620_65240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6663 n_58520_65240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6664 n_59660_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6665 n_66880_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6666 n_63460_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6667 n_63080_65240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6668 n_61940_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6669 n_55100_56840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6670 n_46360_76440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6671 n_40660_76440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6672 n_40660_70840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6673 n_63460_70840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6674 n_74100_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6675 n_65360_70840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6676 n_68780_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6677 n_75240_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6678 n_72960_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6679 n_55480_48440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6680 n_48260_76440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6681 n_45600_84840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6682 n_49400_79240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6683 n_70300_48440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6684 n_40660_79240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6685 n_40280_82040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6686 n_43700_79240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6687 n_44080_84840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6688 n_49400_82040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6689 n_54720_84840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6690 n_44080_59640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6691 n_42940_82040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6692 n_42940_84840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6693 n_40280_84840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6694 n_41420_87640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6695 n_46740_87640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6696 n_43320_87640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6697 n_63080_84840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6698 n_49400_87640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6699 n_64220_82040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6700 n_43320_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6701 n_43320_76440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6702 n_41800_82040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6703 n_68780_56840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6704 n_51680_84840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6705 n_54340_76440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6706 n_65740_82040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6707 n_56240_76440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6708 n_60040_54040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6709 n_68780_59640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6710 n_67260_56840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6711 n_66880_59640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6712 n_70300_59640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6713 n_70300_56840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6714 n_71820_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6715 n_73720_65240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6716 n_70300_70840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6717 n_70300_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6718 n_67260_76440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6719 n_68780_76440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6720 n_59660_82040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6721 n_88920_62440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6722 n_87020_59640 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6723 n_83220_62440 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6724 n_83220_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6725 n_84740_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6726 n_83600_70840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6727 n_85500_70840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6728 n_85880_68040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6729 n_85500_82040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6730 n_68780_82040 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6731 n_43320_65240 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6732 n_44460_56840 0 PWL(54000ps 0uA 54030ps 0uA 54031ps 30uA 54059ps 30uA 54060ps 0uA)
I6733 n_90820_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6734 n_93480_79240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6735 n_91960_87640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6736 n_87020_87640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6737 n_93480_73640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6738 n_93100_84840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6739 n_65740_40040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6740 n_56240_48440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6741 n_40280_54040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6742 n_40660_56840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6743 n_93480_48440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6744 n_92340_48440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6745 n_41800_42840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6746 n_50920_48440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6747 n_70300_40040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6748 n_56620_40040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6749 n_67260_40040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6750 n_93480_45640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6751 n_80560_40040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6752 n_40280_48440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6753 n_72200_40040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6754 n_77140_40040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6755 n_50160_59640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6756 n_42180_73640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6757 n_45600_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6758 n_43320_62440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6759 n_40660_65240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6760 n_41800_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6761 n_44460_62440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6762 n_47500_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6763 n_52060_73640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6764 n_51300_59640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6765 n_74860_40040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6766 n_71820_42840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6767 n_41420_48440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6768 n_80180_42840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6769 n_88920_45640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6770 n_66880_45640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6771 n_57760_40040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6772 n_68400_40040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6773 n_51680_48440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6774 n_48260_45640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6775 n_85120_48440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6776 n_90440_48440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6777 n_41420_54040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6778 n_47880_54040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6779 n_55100_54040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6780 n_63080_51240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6781 n_90820_84840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6782 n_90440_73640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6783 n_85120_84840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6784 n_87400_84840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6785 n_91580_79240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6786 n_88540_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6787 n_87780_54040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6788 n_88920_51240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6789 n_83220_54040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6790 n_91200_54040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6791 n_87400_65240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6792 n_92720_82040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6793 n_88920_82040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6794 n_82080_84840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6795 n_83600_51240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6796 n_80560_51240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6797 n_84740_54040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6798 n_87400_56840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6799 n_90820_56840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6800 n_77520_54040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6801 n_87400_79240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6802 n_88920_65240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6803 n_91960_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6804 n_92340_73640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6805 n_89300_84840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6806 n_81700_82040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6807 n_79040_87640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6808 n_79040_54040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6809 n_80560_54040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6810 n_82080_54040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6811 n_80180_59640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6812 n_76380_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6813 n_67260_84840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6814 n_71820_79240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6815 n_67260_87640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6816 n_65740_84840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6817 n_62320_82040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6818 n_68780_87640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6819 n_71820_87640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6820 n_70300_87640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6821 n_85500_56840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6822 n_85500_59640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6823 n_84740_65240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6824 n_82080_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6825 n_87400_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6826 n_82080_70840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6827 n_77140_70840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6828 n_81700_73640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6829 n_81700_76440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6830 n_72200_76440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6831 n_76760_79240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6832 n_60800_51240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6833 n_53580_54040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6834 n_46360_54040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6835 n_41800_56840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6836 n_87400_51240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6837 n_83600_48440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6838 n_49400_48440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6839 n_53200_48440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6840 n_70300_42840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6841 n_61560_40040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6842 n_68020_48440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6843 n_88920_42840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6844 n_82080_42840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6845 n_42940_48440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6846 n_73720_45640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6847 n_73340_40040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6848 n_57000_54040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6849 n_48260_65240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6850 n_50920_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6851 n_53580_59640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6852 n_53580_62440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6853 n_52060_65240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6854 n_49400_65240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6855 n_56620_65240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6856 n_58520_65240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6857 n_59660_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6858 n_66880_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6859 n_63080_65240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6860 n_61940_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6861 n_55100_56840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6862 n_69160_62440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6863 n_55100_70840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6864 n_53580_70840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6865 n_50920_70840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6866 n_50920_73640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6867 n_49400_73640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6868 n_55860_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6869 n_48260_73640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6870 n_49780_76440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6871 n_50920_79240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6872 n_58520_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6873 n_74100_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6874 n_75240_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6875 n_45600_84840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6876 n_48640_79240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6877 n_60040_76440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6878 n_56620_79240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6879 n_52060_82040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6880 n_70300_48440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6881 n_46360_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6882 n_44840_70840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6883 n_43320_70840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6884 n_41800_70840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6885 n_40660_79240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6886 n_40280_82040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6887 n_44080_84840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6888 n_57380_76440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6889 n_50920_82040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6890 n_50160_84840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6891 n_47500_56840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6892 n_52820_79240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6893 n_44080_59640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6894 n_42940_82040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6895 n_42940_84840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6896 n_40280_84840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6897 n_41420_87640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6898 n_46740_87640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6899 n_43320_87640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6900 n_46740_84840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6901 n_52440_87640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6902 n_59660_84840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6903 n_43320_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6904 n_43320_76440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6905 n_41800_82040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6906 n_51680_84840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6907 n_60800_84840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6908 n_60800_87640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6909 n_74860_87640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6910 n_54340_76440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6911 n_54340_87640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6912 n_64600_84840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6913 n_73340_87640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6914 n_56240_76440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6915 n_71820_59640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6916 n_70300_65240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6917 n_68400_65240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6918 n_71820_65240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6919 n_71820_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6920 n_70300_70840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6921 n_70300_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6922 n_67260_76440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6923 n_65740_79240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6924 n_53960_79240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6925 n_55100_79240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6926 n_59660_82040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6927 n_87020_59640 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6928 n_83220_62440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6929 n_83220_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6930 n_83600_70840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6931 n_85500_70840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6932 n_85880_68040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6933 n_85500_76440 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6934 n_85500_79240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6935 n_83600_82040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6936 n_69920_82040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6937 n_71060_82040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6938 n_72200_82040 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6939 n_43320_65240 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6940 n_44460_56840 0 PWL(56000ps 0uA 56030ps 0uA 56031ps 30uA 56059ps 30uA 56060ps 0uA)
I6941 n_92340_54040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6942 n_93480_62440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6943 n_93480_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6944 n_93100_87640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6945 n_93480_68040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6946 n_93480_73640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6947 n_93100_84840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6948 n_83600_87640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6949 n_65740_40040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6950 n_61940_48440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6951 n_40280_54040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6952 n_44080_54040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6953 n_92340_48440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6954 n_41800_42840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6955 n_48640_40040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6956 n_50920_48440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6957 n_91580_40040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6958 n_52440_40040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6959 n_40660_42840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6960 n_90440_40040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6961 n_80560_40040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6962 n_46360_40040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6963 n_72200_40040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6964 n_82080_48440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6965 n_50160_59640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6966 n_44460_68040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6967 n_45600_68040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6968 n_40660_65240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6969 n_41800_68040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6970 n_47500_68040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6971 n_46740_65240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6972 n_51300_59640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6973 n_80180_45640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6974 n_71820_42840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6975 n_49400_40040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6976 n_80180_42840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6977 n_83600_42840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6978 n_43700_42840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6979 n_51680_42840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6980 n_92720_40040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6981 n_51680_48440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6982 n_47880_42840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6983 n_48260_45640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6984 n_85120_48440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6985 n_49020_51240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6986 n_47880_54040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6987 n_60040_48440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6988 n_63080_51240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6989 n_80180_87640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6990 n_90820_84840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6991 n_90440_73640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6992 n_92340_65240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6993 n_90060_87640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6994 n_91580_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6995 n_91580_62440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6996 n_89300_54040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6997 n_68780_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6998 n_87780_54040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I6999 n_83220_54040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7000 n_91200_54040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7001 n_90820_65240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7002 n_92720_82040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7003 n_85880_87640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7004 n_83600_51240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7005 n_80560_51240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7006 n_84740_54040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7007 n_87400_56840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7008 n_90820_56840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7009 n_77520_54040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7010 n_87400_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7011 n_91960_68040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7012 n_92340_73640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7013 n_89300_84840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7014 n_80560_84840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7015 n_81700_82040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7016 n_79040_87640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7017 n_79040_54040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7018 n_80560_54040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7019 n_82080_54040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7020 n_76380_68040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7021 n_78280_70840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7022 n_75240_76440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7023 n_73720_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7024 n_73720_73640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7025 n_67260_84840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7026 n_71820_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7027 n_88920_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7028 n_67260_87640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7029 n_65740_84840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7030 n_62320_82040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7031 n_68780_87640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7032 n_71820_87640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7033 n_70300_87640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7034 n_70300_84840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7035 n_73720_82040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7036 n_85500_56840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7037 n_86260_54040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7038 n_87400_48440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7039 n_82080_59640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7040 n_82080_65240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7041 n_81700_76440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7042 n_78660_73640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7043 n_78660_76440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7044 n_78660_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7045 n_72200_76440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7046 n_78280_82040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7047 n_76760_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7048 n_80560_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7049 n_80180_82040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7050 n_76760_84840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7051 n_78660_84840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7052 n_74860_82040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7053 n_76760_82040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7054 n_67260_51240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7055 n_71820_51240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7056 n_71820_54040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7057 n_59280_51240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7058 n_49780_54040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7059 n_50920_51240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7060 n_41800_56840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7061 n_52060_51240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7062 n_70300_54040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7063 n_61560_54040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7064 n_83600_48440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7065 n_49400_48440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7066 n_51680_45640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7067 n_53200_48440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7068 n_92720_42840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7069 n_50540_42840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7070 n_45220_42840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7071 n_85500_42840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7072 n_82080_42840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7073 n_51300_40040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7074 n_73720_45640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7075 n_82080_45640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7076 n_48260_65240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7077 n_50920_68040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7078 n_72200_56840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7079 n_53580_59640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7080 n_53580_62440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7081 n_52060_65240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7082 n_49400_65240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7083 n_56620_65240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7084 n_58520_65240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7085 n_60420_65240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7086 n_73720_62440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7087 n_63460_68040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7088 n_60040_73640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7089 n_75240_62440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7090 n_76380_59640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7091 n_63080_82040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7092 n_75240_59640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7093 n_73340_59640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7094 n_61940_68040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7095 n_59660_70840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7096 n_46360_76440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7097 n_48260_73640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7098 n_58520_68040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7099 n_58520_73640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7100 n_56620_73640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7101 n_58140_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7102 n_63460_70840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7103 n_65360_70840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7104 n_68780_68040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7105 n_68020_62440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7106 n_53580_65240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7107 n_53580_68040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7108 n_49400_70840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7109 n_46740_70840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7110 n_48260_76440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7111 n_47500_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7112 n_45600_84840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7113 n_48640_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7114 n_58520_70840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7115 n_60040_76440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7116 n_60420_70840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7117 n_63080_73640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7118 n_71820_73640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7119 n_76760_73640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7120 n_60040_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7121 n_61560_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7122 n_65740_76440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7123 n_58140_51240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7124 n_70300_48440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7125 n_46360_68040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7126 n_44840_70840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7127 n_43320_70840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7128 n_41800_70840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7129 n_40660_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7130 n_40280_82040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7131 n_44080_84840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7132 n_40280_87640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7133 n_57380_76440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7134 n_63080_76440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7135 n_67260_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7136 n_70300_76440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7137 n_43320_87640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7138 n_58140_87640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7139 n_59660_84840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7140 n_55100_82040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7141 n_61940_87640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7142 n_46740_51240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7143 n_43320_68040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7144 n_43320_76440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7145 n_41800_82040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7146 n_66880_62440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7147 n_65360_54040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7148 n_65360_56840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7149 n_63080_54040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7150 n_59280_87640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7151 n_54340_76440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7152 n_53580_87640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7153 n_58520_84840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7154 n_63460_87640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7155 n_67260_65240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7156 n_63460_62440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7157 n_71820_65240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7158 n_71820_68040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7159 n_70300_70840 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7160 n_67260_76440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7161 n_65740_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7162 n_64600_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7163 n_57380_82040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7164 n_55100_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7165 n_58520_82040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7166 n_59660_82040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7167 n_56240_82040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7168 n_88920_62440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7169 n_83220_62440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7170 n_84740_68040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7171 n_85880_73640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7172 n_81700_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7173 n_85500_76440 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7174 n_85500_79240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7175 n_83600_82040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7176 n_85500_82040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7177 n_69920_82040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7178 n_71060_82040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7179 n_72200_82040 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7180 n_43320_65240 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7181 n_60040_59640 0 PWL(58000ps 0uA 58030ps 0uA 58031ps 30uA 58059ps 30uA 58060ps 0uA)
I7182 n_90820_68040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7183 n_91200_70840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7184 n_93480_79240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7185 n_91960_87640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7186 n_87020_87640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7187 n_93480_56840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7188 n_90440_62440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7189 n_93480_68040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7190 n_93480_73640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7191 n_83600_87640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7192 n_65740_40040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7193 n_54720_48440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7194 n_56240_48440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7195 n_65740_45640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7196 n_44080_54040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7197 n_63840_45640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7198 n_79040_42840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7199 n_93480_48440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7200 n_93480_54040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7201 n_48640_40040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7202 n_63840_40040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7203 n_87020_40040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7204 n_88160_40040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7205 n_42940_42840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7206 n_90440_40040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7207 n_93480_45640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7208 n_46360_40040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7209 n_40280_48440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7210 n_72200_40040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7211 n_77140_40040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7212 n_55100_40040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7213 n_40660_51240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7214 n_44460_68040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7215 n_45600_68040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7216 n_43320_62440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7217 n_44460_62440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7218 n_47500_68040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7219 n_46740_65240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7220 n_44840_51240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7221 n_54720_42840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7222 n_74860_40040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7223 n_71820_42840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7224 n_41420_48440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7225 n_49400_40040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7226 n_88920_45640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7227 n_83600_42840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7228 n_44840_45640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7229 n_83600_40040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7230 n_87020_45640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7231 n_63460_42840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7232 n_47880_42840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7233 n_92340_51240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7234 n_90440_48440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7235 n_78280_48440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7236 n_64980_48440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7237 n_49020_51240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7238 n_64600_51240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7239 n_55100_54040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7240 n_54720_51240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7241 n_63080_51240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7242 n_80180_87640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7243 n_90440_73640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7244 n_92340_65240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7245 n_90820_59640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7246 n_88920_56840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7247 n_85120_84840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7248 n_87400_84840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7249 n_91580_79240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7250 n_87400_73640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7251 n_88540_68040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7252 n_87400_65240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7253 n_87400_76440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7254 n_92340_76440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7255 n_88920_82040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7256 n_82080_84840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7257 n_87400_56840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7258 n_89300_59640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7259 n_88920_65240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7260 n_89300_73640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7261 n_80560_84840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7262 n_76380_54040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7263 n_76760_56840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7264 n_78280_70840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7265 n_73720_70840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7266 n_75240_76440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7267 n_73720_79240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7268 n_70300_79240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7269 n_67260_84840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7270 n_88920_79240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7271 n_67260_87640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7272 n_65740_84840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7273 n_65360_87640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7274 n_70300_84840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7275 n_73720_82040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7276 n_72200_84840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7277 n_86260_54040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7278 n_84740_65240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7279 n_82080_68040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7280 n_87400_68040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7281 n_82080_70840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7282 n_77140_70840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7283 n_81700_73640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7284 n_80560_73640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7285 n_78660_73640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7286 n_78660_76440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7287 n_78660_79240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7288 n_76760_76440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7289 n_78280_82040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7290 n_80560_79240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7291 n_80180_82040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7292 n_76760_84840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7293 n_78660_84840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7294 n_74860_82040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7295 n_76760_82040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7296 n_67260_51240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7297 n_70300_51240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7298 n_68020_54040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7299 n_68780_51240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7300 n_50920_51240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7301 n_66120_51240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7302 n_79040_51240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7303 n_87400_51240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7304 n_90820_51240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7305 n_51680_45640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7306 n_65360_42840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7307 n_90440_45640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7308 n_85500_40040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7309 n_46740_45640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7310 n_85500_42840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7311 n_88920_42840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7312 n_51300_40040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7313 n_42940_48440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7314 n_73720_45640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7315 n_73340_40040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7316 n_53200_42840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7317 n_43320_51240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7318 n_58900_48440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7319 n_72200_56840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7320 n_63460_68040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7321 n_60040_73640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7322 n_75240_59640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7323 n_77520_62440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7324 n_72200_62440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7325 n_61940_68040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7326 n_59660_70840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7327 n_46360_76440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7328 n_48260_73640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7329 n_58520_68040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7330 n_61560_73640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7331 n_70300_73640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7332 n_56620_73640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7333 n_66880_73640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7334 n_58140_79240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7335 n_74100_68040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7336 n_75240_65240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7337 n_55480_48440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7338 n_68780_70840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7339 n_53580_65240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7340 n_53580_68040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7341 n_49400_70840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7342 n_46740_70840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7343 n_48260_76440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7344 n_47500_79240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7345 n_48640_79240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7346 n_58520_70840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7347 n_60040_76440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7348 n_60420_70840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7349 n_71820_73640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7350 n_60040_79240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7351 n_61560_79240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7352 n_52060_82040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7353 n_67260_70840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7354 n_46360_68040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7355 n_44840_70840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7356 n_43320_70840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7357 n_41800_70840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7358 n_40660_79240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7359 n_43700_79240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7360 n_40280_87640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7361 n_57380_76440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7362 n_80560_76440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7363 n_50920_82040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7364 n_50160_84840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7365 n_47500_56840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7366 n_44080_59640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7367 n_42940_82040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7368 n_42940_84840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7369 n_40280_84840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7370 n_41420_87640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7371 n_46740_87640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7372 n_46740_84840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7373 n_52440_87640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7374 n_49400_87640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7375 n_64220_82040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7376 n_58140_87640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7377 n_46740_51240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7378 n_54340_87640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7379 n_67260_82040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7380 n_53580_87640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7381 n_73340_87640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7382 n_57000_87640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7383 n_66880_59640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7384 n_71820_59640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7385 n_68400_65240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7386 n_71820_65240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7387 n_71820_68040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7388 n_70300_70840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7389 n_67260_76440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7390 n_65740_79240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7391 n_64600_79240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7392 n_57380_82040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7393 n_58520_82040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7394 n_59660_82040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7395 n_56240_82040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7396 n_87400_62440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7397 n_87020_59640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7398 n_88160_59640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7399 n_85880_62440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7400 n_83220_65240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7401 n_84740_62440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7402 n_83220_68040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7403 n_84740_68040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7404 n_83600_70840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7405 n_85500_70840 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7406 n_83220_73640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7407 n_84740_73640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7408 n_85880_68040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7409 n_85880_73640 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7410 n_83600_76440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7411 n_85500_76440 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7412 n_85500_79240 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7413 n_87400_82040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7414 n_83600_82040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7415 n_85500_82040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7416 n_69920_82040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7417 n_71060_82040 0 PWL(60000ps 0uA 60030ps 0uA 60031ps 30uA 60059ps 30uA 60060ps 0uA)
I7418 n_92340_54040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7419 n_93480_62440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7420 n_90820_68040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7421 n_93480_79240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7422 n_93100_87640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7423 n_93480_56840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7424 n_93480_73640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7425 n_93480_76440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7426 n_83600_87640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7427 n_84740_87640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7428 n_65740_40040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7429 n_54720_48440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7430 n_56240_48440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7431 n_44080_54040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7432 n_40660_56840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7433 n_63840_45640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7434 n_79040_42840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7435 n_93480_48440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7436 n_48640_40040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7437 n_50920_48440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7438 n_63840_40040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7439 n_52440_40040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7440 n_40660_42840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7441 n_56620_40040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7442 n_67260_40040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7443 n_90440_40040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7444 n_93480_45640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7445 n_40280_40040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7446 n_82080_48440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7447 n_55100_40040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7448 n_40660_51240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7449 n_44460_68040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7450 n_45600_68040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7451 n_43320_62440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7452 n_40660_65240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7453 n_41800_68040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7454 n_44460_62440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7455 n_47500_68040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7456 n_46740_65240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7457 n_44840_51240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7458 n_54720_42840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7459 n_80180_45640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7460 n_41420_40040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7461 n_88920_45640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7462 n_83600_42840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7463 n_66880_45640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7464 n_57760_40040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7465 n_43700_42840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7466 n_51680_42840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7467 n_63460_42840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7468 n_51680_48440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7469 n_47880_42840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7470 n_90440_48440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7471 n_78280_48440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7472 n_64980_48440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7473 n_41420_54040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7474 n_49020_51240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7475 n_55100_54040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7476 n_54720_51240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7477 n_63080_51240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7478 n_81700_87640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7479 n_80180_87640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7480 n_90440_76440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7481 n_90440_73640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7482 n_88920_56840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7483 n_90060_87640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7484 n_91580_79240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7485 n_88540_68040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7486 n_91580_62440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7487 n_89300_54040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7488 n_87780_54040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7489 n_83220_54040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7490 n_91200_54040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7491 n_90820_65240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7492 n_87400_65240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7493 n_87400_70840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7494 n_87400_76440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7495 n_92340_76440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7496 n_87780_87640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7497 n_88920_82040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7498 n_83600_84840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7499 n_82080_84840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7500 n_85880_87640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7501 n_83600_51240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7502 n_80560_51240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7503 n_84740_54040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7504 n_90820_56840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7505 n_77520_54040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7506 n_87400_79240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7507 n_89300_59640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7508 n_92720_59640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7509 n_88920_65240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7510 n_91960_68040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7511 n_89300_73640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7512 n_90060_79240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7513 n_89300_84840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7514 n_90820_82040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7515 n_77900_87640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7516 n_81700_82040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7517 n_79040_54040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7518 n_80560_54040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7519 n_82080_54040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7520 n_76380_54040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7521 n_76760_56840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7522 n_76380_68040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7523 n_80560_65240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7524 n_77900_68040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7525 n_76000_70840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7526 n_74860_70840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7527 n_75240_76440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7528 n_73720_79240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7529 n_70300_79240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7530 n_67260_84840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7531 n_88920_79240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7532 n_67260_87640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7533 n_65360_87640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7534 n_70300_87640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7535 n_73720_82040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7536 n_85500_56840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7537 n_87400_48440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7538 n_82080_59640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7539 n_84740_65240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7540 n_82080_65240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7541 n_82080_68040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7542 n_87400_68040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7543 n_82080_70840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7544 n_77140_70840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7545 n_81700_73640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7546 n_78660_73640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7547 n_78660_76440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7548 n_78660_79240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7549 n_76760_76440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7550 n_78280_82040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7551 n_80560_79240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7552 n_76760_84840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7553 n_78660_84840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7554 n_74860_82040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7555 n_67260_51240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7556 n_70300_51240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7557 n_68020_54040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7558 n_50920_51240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7559 n_52060_51240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7560 n_66120_51240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7561 n_79040_51240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7562 n_87400_51240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7563 n_51680_45640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7564 n_53200_48440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7565 n_65360_42840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7566 n_50540_42840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7567 n_45220_42840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7568 n_61560_40040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7569 n_68020_48440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7570 n_85500_42840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7571 n_88920_42840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7572 n_43320_40040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7573 n_82080_45640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7574 n_53200_42840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7575 n_43320_51240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7576 n_58900_48440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7577 n_57000_54040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7578 n_52060_54040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7579 n_72200_56840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7580 n_63460_68040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7581 n_75240_59640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7582 n_72200_62440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7583 n_55100_56840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7584 n_55860_68040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7585 n_46740_73640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7586 n_40660_76440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7587 n_48260_73640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7588 n_40660_70840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7589 n_49780_76440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7590 n_50920_79240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7591 n_58520_68040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7592 n_74100_68040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7593 n_75240_65240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7594 n_55480_48440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7595 n_53580_65240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7596 n_53580_68040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7597 n_49400_70840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7598 n_46740_70840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7599 n_46360_68040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7600 n_44840_70840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7601 n_43320_70840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7602 n_41800_70840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7603 n_40280_82040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7604 n_44080_84840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7605 n_80560_76440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7606 n_47500_56840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7607 n_44080_59640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7608 n_42940_82040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7609 n_42940_84840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7610 n_40280_84840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7611 n_49400_87640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7612 n_64220_82040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7613 n_43320_68040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7614 n_43320_76440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7615 n_41800_82040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7616 n_45220_87640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7617 n_51680_84840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7618 n_67260_82040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7619 n_66880_59640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7620 n_71820_59640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7621 n_68400_65240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7622 n_59660_82040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7623 n_87400_62440 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7624 n_87020_59640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7625 n_88160_59640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7626 n_83220_65240 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7627 n_83220_73640 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7628 n_85880_68040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7629 n_87400_82040 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7630 n_44460_56840 0 PWL(62000ps 0uA 62030ps 0uA 62031ps 30uA 62059ps 30uA 62060ps 0uA)
I7631 n_92340_54040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7632 n_93480_62440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7633 n_91200_70840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7634 n_93480_79240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7635 n_93480_56840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7636 n_90440_62440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7637 n_93480_76440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7638 n_83600_87640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7639 n_65740_40040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7640 n_56240_48440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7641 n_65740_45640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7642 n_44080_54040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7643 n_40660_56840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7644 n_63840_45640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7645 n_93480_48440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7646 n_93480_54040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7647 n_48640_40040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7648 n_50920_48440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7649 n_70300_40040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7650 n_91580_40040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7651 n_88160_40040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7652 n_52440_40040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7653 n_40660_42840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7654 n_56620_40040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7655 n_90440_40040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7656 n_93480_45640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7657 n_80560_40040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7658 n_40280_40040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7659 n_40280_48440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7660 n_60040_45640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7661 n_72200_40040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7662 n_55100_40040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7663 n_54720_42840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7664 n_71820_42840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7665 n_56620_45640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7666 n_41420_48440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7667 n_41420_40040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7668 n_80180_42840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7669 n_88920_45640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7670 n_83600_42840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7671 n_57760_40040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7672 n_43700_42840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7673 n_51680_42840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7674 n_83600_40040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7675 n_92720_40040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7676 n_68400_40040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7677 n_51680_48440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7678 n_47880_42840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7679 n_92340_51240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7680 n_90440_48440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7681 n_64980_48440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7682 n_41420_54040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7683 n_49020_51240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7684 n_64600_51240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7685 n_55100_54040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7686 n_63080_51240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7687 n_80180_87640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7688 n_90440_76440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7689 n_90820_59640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7690 n_88920_56840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7691 n_91580_79240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7692 n_87400_73640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7693 n_91580_62440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7694 n_89300_54040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7695 n_87780_54040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7696 n_83220_54040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7697 n_91200_54040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7698 n_90820_65240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7699 n_87400_70840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7700 n_92340_76440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7701 n_87780_87640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7702 n_88920_82040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7703 n_83600_84840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7704 n_82080_84840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7705 n_83600_51240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7706 n_80560_51240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7707 n_84740_54040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7708 n_90820_56840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7709 n_92720_59640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7710 n_90060_79240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7711 n_77900_87640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7712 n_82080_54040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7713 n_80560_56840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7714 n_82080_56840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7715 n_78660_56840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7716 n_76380_54040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7717 n_76760_65240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7718 n_76380_68040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7719 n_78660_65240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7720 n_80560_65240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7721 n_75240_73640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7722 n_74860_70840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7723 n_73720_70840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7724 n_75240_76440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7725 n_88920_79240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7726 n_70300_87640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7727 n_73720_82040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7728 n_72200_84840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7729 n_85500_56840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7730 n_87400_48440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7731 n_82080_59640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7732 n_82080_65240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7733 n_82080_68040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7734 n_85880_65240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7735 n_82080_70840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7736 n_77140_70840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7737 n_81700_73640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7738 n_80560_73640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7739 n_78660_73640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7740 n_78660_76440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7741 n_78660_79240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7742 n_76760_76440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7743 n_78280_82040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7744 n_80560_79240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7745 n_76760_84840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7746 n_78660_84840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7747 n_74860_82040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7748 n_67260_51240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7749 n_68020_54040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7750 n_68780_51240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7751 n_50920_51240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7752 n_52060_51240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7753 n_66120_51240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7754 n_87400_51240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7755 n_90820_51240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7756 n_51680_45640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7757 n_53200_48440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7758 n_70300_42840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7759 n_92720_42840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7760 n_85500_40040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7761 n_50540_42840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7762 n_45220_42840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7763 n_61560_40040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7764 n_85500_42840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7765 n_88920_42840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7766 n_82080_42840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7767 n_43320_40040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7768 n_42940_48440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7769 n_53200_45640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7770 n_73720_45640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7771 n_53200_42840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7772 n_58900_48440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7773 n_52060_54040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7774 n_72200_56840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7775 n_59660_68040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7776 n_60420_65240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7777 n_73720_62440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7778 n_66880_68040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7779 n_60800_68040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7780 n_63460_68040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7781 n_60040_73640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7782 n_63080_65240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7783 n_75240_62440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7784 n_76380_59640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7785 n_75240_59640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7786 n_72200_62440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7787 n_61940_68040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7788 n_59660_70840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7789 n_55100_56840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7790 n_69160_62440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7791 n_55860_68040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7792 n_46360_79240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7793 n_61560_73640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7794 n_70300_73640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7795 n_56620_73640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7796 n_66880_73640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7797 n_58140_79240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7798 n_63460_70840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7799 n_74100_68040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7800 n_65360_68040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7801 n_68780_68040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7802 n_75240_65240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7803 n_68020_62440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7804 n_55480_48440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7805 n_68780_70840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7806 n_48260_76440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7807 n_47500_79240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7808 n_45600_84840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7809 n_48640_79240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7810 n_58520_70840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7811 n_49400_79240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7812 n_60040_76440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7813 n_60420_70840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7814 n_71820_73640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7815 n_60040_79240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7816 n_61560_79240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7817 n_52060_82040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7818 n_67260_70840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7819 n_58140_51240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7820 n_57380_76440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7821 n_80560_76440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7822 n_50920_82040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7823 n_50160_84840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7824 n_41420_87640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7825 n_46740_87640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7826 n_43320_87640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7827 n_46740_84840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7828 n_52440_87640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7829 n_64220_82040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7830 n_50920_87640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7831 n_58140_87640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7832 n_59660_84840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7833 n_46740_51240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7834 n_45220_87640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7835 n_59280_87640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7836 n_51680_84840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7837 n_74860_87640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7838 n_67260_82040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7839 n_53580_87640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7840 n_58520_84840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7841 n_56240_76440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7842 n_57000_87640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7843 n_66880_59640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7844 n_71820_59640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7845 n_70300_65240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7846 n_68400_65240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7847 n_71820_65240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7848 n_71820_68040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7849 n_70300_70840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7850 n_70300_68040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7851 n_67260_76440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7852 n_65740_79240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7853 n_64600_79240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7854 n_57380_82040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7855 n_58520_82040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7856 n_56240_82040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7857 n_87400_62440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7858 n_87020_59640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7859 n_85880_62440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7860 n_84740_62440 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7861 n_83220_68040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7862 n_83600_70840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7863 n_85500_70840 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7864 n_84740_73640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7865 n_85880_73640 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7866 n_85500_79240 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7867 n_87400_82040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7868 n_83600_82040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7869 n_69920_82040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7870 n_71060_82040 0 PWL(64000ps 0uA 64030ps 0uA 64031ps 30uA 64059ps 30uA 64060ps 0uA)
I7871 n_93480_79240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7872 n_91960_87640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7873 n_93100_87640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7874 n_90440_62440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7875 n_93480_68040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7876 n_93100_84840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7877 n_54720_48440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7878 n_56240_48440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7879 n_40280_54040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7880 n_40660_56840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7881 n_79040_42840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7882 n_93480_48440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7883 n_41800_42840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7884 n_50920_48440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7885 n_63840_40040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7886 n_70300_40040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7887 n_91580_40040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7888 n_87020_40040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7889 n_88160_40040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7890 n_52440_40040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7891 n_40660_42840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7892 n_90440_40040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7893 n_93480_45640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7894 n_46360_40040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7895 n_40280_40040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7896 n_40280_48440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7897 n_72200_40040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7898 n_79040_40040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7899 n_82080_48440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7900 n_43320_59640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7901 n_50160_59640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7902 n_42180_73640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7903 n_52060_73640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7904 n_51300_59640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7905 n_46740_59640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7906 n_80180_45640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7907 n_76760_42840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7908 n_71820_42840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7909 n_41420_48440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7910 n_41420_40040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7911 n_49400_40040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7912 n_88920_45640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7913 n_83600_42840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7914 n_43700_42840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7915 n_51680_42840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7916 n_83600_40040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7917 n_87020_45640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7918 n_92720_40040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7919 n_68400_40040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7920 n_63460_42840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7921 n_51680_48440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7922 n_48260_45640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7923 n_90440_48440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7924 n_78280_48440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7925 n_41420_54040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7926 n_47880_54040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7927 n_55100_54040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7928 n_54720_51240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7929 n_90820_84840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7930 n_92340_65240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7931 n_90820_59640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7932 n_90060_87640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7933 n_87400_84840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7934 n_91580_79240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7935 n_92340_76440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7936 n_88920_82040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7937 n_85880_87640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7938 n_77520_54040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7939 n_87400_79240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7940 n_89300_59640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7941 n_91960_68040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7942 n_90820_82040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7943 n_79040_54040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7944 n_80560_54040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7945 n_80560_56840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7946 n_82080_56840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7947 n_78660_56840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7948 n_76760_65240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7949 n_76760_56840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7950 n_78660_65240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7951 n_77900_68040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7952 n_76000_70840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7953 n_78280_70840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7954 n_75240_73640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7955 n_73720_79240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7956 n_70300_79240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7957 n_67260_84840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7958 n_67260_87640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7959 n_62320_82040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7960 n_68780_87640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7961 n_71820_87640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7962 n_70300_87640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7963 n_84740_65240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7964 n_85880_65240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7965 n_77140_70840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7966 n_76760_76440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7967 n_80560_79240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7968 n_70300_51240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7969 n_68020_54040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7970 n_49780_54040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7971 n_52060_51240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7972 n_79040_51240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7973 n_87400_51240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7974 n_49400_48440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7975 n_53200_48440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7976 n_65360_42840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7977 n_70300_42840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7978 n_92720_42840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7979 n_90440_45640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7980 n_85500_40040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7981 n_50540_42840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7982 n_45220_42840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7983 n_85500_42840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7984 n_88920_42840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7985 n_51300_40040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7986 n_43320_40040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7987 n_42940_48440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7988 n_73720_45640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7989 n_76760_45640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7990 n_82080_45640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7991 n_49780_56840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7992 n_48260_62440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7993 n_49780_62440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7994 n_44840_73640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7995 n_53580_59640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7996 n_53580_62440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7997 n_52060_65240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7998 n_49400_65240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I7999 n_59660_68040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8000 n_60420_65240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8001 n_73720_62440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8002 n_66880_68040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8003 n_60800_68040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8004 n_60040_73640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8005 n_63080_65240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8006 n_75240_62440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8007 n_76380_59640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8008 n_61940_68040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8009 n_59660_70840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8010 n_55100_56840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8011 n_55100_70840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8012 n_53580_70840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8013 n_50920_70840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8014 n_50920_73640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8015 n_48260_73640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8016 n_49780_76440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8017 n_50920_79240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8018 n_46360_79240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8019 n_58520_68040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8020 n_58520_73640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8021 n_56620_73640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8022 n_58140_79240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8023 n_74100_68040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8024 n_75240_65240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8025 n_48260_76440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8026 n_47500_79240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8027 n_45600_84840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8028 n_48640_79240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8029 n_58520_70840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8030 n_49400_79240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8031 n_60040_76440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8032 n_60420_70840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8033 n_63080_73640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8034 n_60040_79240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8035 n_61560_79240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8036 n_52060_82040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8037 n_57380_76440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8038 n_80560_76440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8039 n_49400_82040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8040 n_54720_84840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8041 n_53580_82040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8042 n_50160_84840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8043 n_52820_79240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8044 n_41420_87640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8045 n_46740_87640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8046 n_43320_87640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8047 n_61940_84840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8048 n_49400_84840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8049 n_49400_87640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8050 n_50920_87640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8051 n_59660_84840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8052 n_55100_82040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8053 n_45220_87640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8054 n_59280_87640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8055 n_51680_84840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8056 n_74860_87640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8057 n_54340_87640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8058 n_58520_84840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8059 n_73340_87640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8060 n_56240_76440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8061 n_70300_65240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8062 n_71820_65240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8063 n_71820_68040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8064 n_70300_70840 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8065 n_70300_68040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8066 n_67260_76440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8067 n_65740_79240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8068 n_64600_79240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8069 n_57380_82040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8070 n_58520_82040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8071 n_59660_82040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8072 n_88160_59640 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8073 n_85880_62440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8074 n_84740_62440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8075 n_84740_68040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8076 n_83600_76440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8077 n_81700_79240 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8078 n_85500_76440 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8079 n_87400_82040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8080 n_85500_82040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8081 n_69920_82040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8082 n_71060_82040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8083 n_72200_82040 0 PWL(66000ps 0uA 66030ps 0uA 66031ps 30uA 66059ps 30uA 66060ps 0uA)
I8084 n_93480_62440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8085 n_90820_68040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8086 n_91200_70840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8087 n_93480_79240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8088 n_87020_87640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8089 n_93480_56840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8090 n_90440_62440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8091 n_93480_73640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8092 n_83600_87640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8093 n_65740_40040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8094 n_54720_48440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8095 n_65740_45640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8096 n_40280_54040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8097 n_40660_56840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8098 n_63840_45640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8099 n_79040_42840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8100 n_93480_54040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8101 n_41800_42840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8102 n_50920_48440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8103 n_91580_40040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8104 n_87020_40040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8105 n_52440_40040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8106 n_40660_42840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8107 n_42940_42840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8108 n_56620_40040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8109 n_93480_45640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8110 n_80560_40040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8111 n_40280_40040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8112 n_40280_48440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8113 n_60040_45640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8114 n_72200_40040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8115 n_40660_45640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8116 n_43320_59640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8117 n_42180_73640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8118 n_45600_68040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8119 n_43320_62440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8120 n_44460_62440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8121 n_47500_68040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8122 n_52060_73640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8123 n_46740_59640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8124 n_45220_48440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8125 n_71820_42840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8126 n_56620_45640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8127 n_41420_48440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8128 n_41420_40040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8129 n_80180_42840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8130 n_88920_45640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8131 n_57760_40040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8132 n_44840_45640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8133 n_43700_42840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8134 n_51680_42840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8135 n_87020_45640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8136 n_92720_40040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8137 n_51680_48440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8138 n_48260_45640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8139 n_92340_51240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8140 n_78280_48440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8141 n_64980_48440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8142 n_41420_54040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8143 n_47880_54040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8144 n_64600_51240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8145 n_54720_51240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8146 n_63080_51240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8147 n_80180_87640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8148 n_90440_73640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8149 n_90820_59640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8150 n_88920_56840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8151 n_85120_84840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8152 n_91580_79240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8153 n_87400_73640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8154 n_88540_68040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8155 n_91580_62440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8156 n_90820_65240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8157 n_87400_65240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8158 n_87400_76440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8159 n_92340_76440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8160 n_82080_84840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8161 n_90820_56840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8162 n_77520_54040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8163 n_87400_79240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8164 n_89300_59640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8165 n_92340_73640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8166 n_77900_87640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8167 n_79040_54040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8168 n_80560_54040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8169 n_80560_56840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8170 n_82080_56840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8171 n_78660_56840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8172 n_76380_54040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8173 n_76760_65240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8174 n_76760_56840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8175 n_78660_65240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8176 n_77900_68040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8177 n_76000_70840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8178 n_75240_73640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8179 n_73720_70840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8180 n_73720_79240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8181 n_70300_79240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8182 n_67260_84840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8183 n_65740_84840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8184 n_62320_82040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8185 n_65360_87640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8186 n_68780_87640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8187 n_71820_87640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8188 n_70300_87640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8189 n_72200_84840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8190 n_86260_54040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8191 n_82080_59640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8192 n_85500_59640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8193 n_82080_65240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8194 n_87400_68040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8195 n_80560_68040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8196 n_80560_73640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8197 n_78660_79240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8198 n_76760_76440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8199 n_78280_82040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8200 n_76760_84840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8201 n_78660_84840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8202 n_74860_82040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8203 n_76760_82040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8204 n_67260_51240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8205 n_70300_51240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8206 n_68780_51240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8207 n_49780_54040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8208 n_52060_51240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8209 n_66120_51240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8210 n_79040_51240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8211 n_90820_51240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8212 n_49400_48440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8213 n_53200_48440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8214 n_92720_42840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8215 n_90440_45640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8216 n_50540_42840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8217 n_45220_42840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8218 n_46740_45640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8219 n_61560_40040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8220 n_88920_42840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8221 n_82080_42840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8222 n_43320_40040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8223 n_42940_48440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8224 n_53200_45640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8225 n_73720_45640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8226 n_44080_48440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8227 n_58900_48440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8228 n_57000_54040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8229 n_49780_56840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8230 n_48260_62440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8231 n_48260_65240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8232 n_49780_62440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8233 n_44840_73640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8234 n_50920_68040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8235 n_56620_65240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8236 n_58520_65240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8237 n_60420_65240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8238 n_73720_62440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8239 n_63460_68040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8240 n_60040_73640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8241 n_75240_62440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8242 n_76380_59640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8243 n_77520_62440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8244 n_61940_68040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8245 n_59660_70840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8246 n_69160_62440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8247 n_55100_70840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8248 n_53580_70840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8249 n_50920_70840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8250 n_50920_73640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8251 n_46740_73640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8252 n_46360_76440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8253 n_40660_76440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8254 n_48260_73640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8255 n_40660_70840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8256 n_58520_68040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8257 n_58520_73640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8258 n_70300_73640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8259 n_63460_70840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8260 n_65360_68040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8261 n_68780_68040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8262 n_68020_62440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8263 n_55480_48440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8264 n_48260_76440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8265 n_58520_70840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8266 n_60420_70840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8267 n_71820_73640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8268 n_52060_82040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8269 n_65740_76440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8270 n_58140_51240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8271 n_70300_48440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8272 n_46360_68040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8273 n_44840_70840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8274 n_43320_70840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8275 n_41800_70840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8276 n_40280_82040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8277 n_40280_87640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8278 n_80560_76440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8279 n_49400_82040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8280 n_54720_84840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8281 n_47120_82040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8282 n_50160_84840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8283 n_65740_73640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8284 n_44080_59640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8285 n_42940_82040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8286 n_42940_84840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8287 n_40280_84840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8288 n_41420_87640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8289 n_43320_87640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8290 n_46740_84840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8291 n_61940_84840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8292 n_49400_87640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8293 n_50920_87640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8294 n_59660_84840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8295 n_42940_54040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8296 n_45220_87640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8297 n_59280_87640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8298 n_51680_84840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8299 n_54340_87640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8300 n_58520_84840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8301 n_73340_87640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8302 n_56240_76440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8303 n_66880_59640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8304 n_71820_59640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8305 n_68400_65240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8306 n_71820_65240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8307 n_73720_65240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8308 n_68780_76440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8309 n_65740_79240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8310 n_64600_79240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8311 n_53960_79240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8312 n_57380_82040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8313 n_58520_82040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8314 n_59660_82040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8315 n_87400_62440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8316 n_87020_59640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8317 n_88160_59640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8318 n_85880_62440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8319 n_84740_62440 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8320 n_83220_68040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8321 n_84740_68040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8322 n_83600_70840 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8323 n_83220_73640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8324 n_85880_73640 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8325 n_81700_79240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8326 n_69920_82040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8327 n_68780_82040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8328 n_72200_82040 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8329 n_43320_65240 0 PWL(68000ps 0uA 68030ps 0uA 68031ps 30uA 68059ps 30uA 68060ps 0uA)
I8330 n_93480_62440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8331 n_90820_68040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8332 n_91200_70840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8333 n_87020_87640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8334 n_93100_87640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8335 n_93480_68040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8336 n_93480_73640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8337 n_93480_76440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8338 n_56240_48440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8339 n_65740_45640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8340 n_61940_48440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8341 n_40280_54040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8342 n_44080_54040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8343 n_40660_56840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8344 n_93480_48440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8345 n_93480_54040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8346 n_92340_48440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8347 n_41800_42840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8348 n_48640_40040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8349 n_50920_48440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8350 n_63840_40040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8351 n_91580_40040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8352 n_56620_40040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8353 n_67260_40040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8354 n_90440_40040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8355 n_93480_45640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8356 n_80560_40040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8357 n_46360_40040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8358 n_40280_48440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8359 n_79040_40040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8360 n_40660_45640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8361 n_40660_51240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8362 n_43320_59640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8363 n_42180_73640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8364 n_45600_68040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8365 n_43320_62440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8366 n_44460_62440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8367 n_47500_68040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8368 n_52060_73640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8369 n_46740_59640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8370 n_44840_51240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8371 n_45220_48440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8372 n_76760_42840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8373 n_41420_48440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8374 n_49400_40040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8375 n_80180_42840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8376 n_88920_45640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8377 n_83600_42840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8378 n_66880_45640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8379 n_57760_40040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8380 n_92720_40040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8381 n_63460_42840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8382 n_51680_48440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8383 n_47880_42840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8384 n_48260_45640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8385 n_85120_48440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8386 n_92340_51240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8387 n_90440_48440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8388 n_41420_54040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8389 n_49020_51240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8390 n_47880_54040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8391 n_60040_48440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8392 n_64600_51240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8393 n_55100_54040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8394 n_90440_76440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8395 n_90440_73640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8396 n_92340_65240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8397 n_90060_87640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8398 n_85120_84840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8399 n_87400_73640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8400 n_88540_68040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8401 n_91580_62440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8402 n_68780_79240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8403 n_90820_65240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8404 n_87400_65240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8405 n_87400_76440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8406 n_82080_84840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8407 n_85880_87640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8408 n_87400_56840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8409 n_90820_56840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8410 n_77520_54040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8411 n_87400_79240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8412 n_88920_65240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8413 n_92340_73640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8414 n_88920_76440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8415 n_80560_84840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8416 n_77900_87640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8417 n_79040_54040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8418 n_80560_54040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8419 n_80560_56840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8420 n_82080_56840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8421 n_78660_56840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8422 n_76760_65240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8423 n_78660_65240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8424 n_77900_68040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8425 n_76000_70840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8426 n_78280_70840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8427 n_75240_73640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8428 n_73720_70840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8429 n_73720_79240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8430 n_73720_73640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8431 n_67260_84840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8432 n_71820_79240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8433 n_65740_84840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8434 n_62320_82040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8435 n_65360_87640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8436 n_68780_87640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8437 n_68780_84840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8438 n_70300_84840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8439 n_73720_82040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8440 n_72200_84840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8441 n_82080_59640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8442 n_85500_59640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8443 n_84740_65240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8444 n_82080_65240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8445 n_85880_65240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8446 n_87400_68040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8447 n_80560_68040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8448 n_77140_70840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8449 n_80560_73640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8450 n_78660_79240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8451 n_76760_76440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8452 n_72200_76440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8453 n_78280_82040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8454 n_76760_84840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8455 n_78660_84840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8456 n_74860_84840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8457 n_76760_82040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8458 n_68020_54040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8459 n_68780_51240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8460 n_61940_51240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8461 n_49780_54040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8462 n_50920_51240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8463 n_52060_51240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8464 n_87400_51240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8465 n_90820_51240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8466 n_83600_48440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8467 n_49400_48440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8468 n_51680_45640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8469 n_53200_48440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8470 n_65360_42840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8471 n_92720_42840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8472 n_61560_40040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8473 n_68020_48440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8474 n_85500_42840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8475 n_88920_42840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8476 n_82080_42840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8477 n_51300_40040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8478 n_42940_48440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8479 n_76760_45640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8480 n_44080_48440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8481 n_43320_51240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8482 n_49780_56840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8483 n_48260_62440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8484 n_48260_65240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8485 n_49780_62440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8486 n_44840_73640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8487 n_50920_68040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8488 n_56620_65240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8489 n_58520_65240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8490 n_60420_65240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8491 n_73720_62440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8492 n_63460_68040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8493 n_60040_73640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8494 n_76380_62440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8495 n_63080_82040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8496 n_77520_62440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8497 n_72200_62440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8498 n_73340_59640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8499 n_61940_68040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8500 n_59660_70840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8501 n_55100_56840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8502 n_55100_70840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8503 n_53580_70840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8504 n_50920_70840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8505 n_50920_73640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8506 n_46740_73640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8507 n_46360_76440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8508 n_40660_76440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8509 n_48260_73640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8510 n_40660_70840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8511 n_58520_68040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8512 n_58520_73640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8513 n_70300_73640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8514 n_63460_70840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8515 n_65360_70840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8516 n_68780_68040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8517 n_68020_62440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8518 n_55480_48440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8519 n_48260_76440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8520 n_58520_70840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8521 n_60420_70840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8522 n_76760_73640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8523 n_56620_79240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8524 n_60040_79240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8525 n_63080_79240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8526 n_52060_82040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8527 n_46360_68040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8528 n_44840_70840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8529 n_43320_70840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8530 n_41800_70840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8531 n_40280_82040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8532 n_40280_87640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8533 n_57380_76440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8534 n_63080_76440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8535 n_49400_82040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8536 n_54720_84840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8537 n_47120_82040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8538 n_50160_84840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8539 n_65740_73640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8540 n_70300_76440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8541 n_52820_79240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8542 n_44080_59640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8543 n_42940_82040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8544 n_42940_84840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8545 n_40280_84840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8546 n_41420_87640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8547 n_43320_87640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8548 n_46740_84840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8549 n_63080_84840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8550 n_52440_87640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8551 n_64220_82040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8552 n_50920_87640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8553 n_58140_87640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8554 n_59660_84840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8555 n_42940_54040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8556 n_46740_51240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8557 n_66880_62440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8558 n_65360_54040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8559 n_63080_54040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8560 n_45220_87640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8561 n_59280_87640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8562 n_51680_84840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8563 n_67260_82040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8564 n_53580_87640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8565 n_64600_84840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8566 n_56240_76440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8567 n_63460_87640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8568 n_67260_65240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8569 n_63460_62440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8570 n_60040_54040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8571 n_68400_65240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8572 n_71820_65240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8573 n_73720_65240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8574 n_68780_76440 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8575 n_65740_79240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8576 n_64600_79240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8577 n_53960_79240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8578 n_57380_82040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8579 n_55100_79240 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8580 n_58520_82040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8581 n_56240_82040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8582 n_83220_68040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8583 n_83600_70840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8584 n_83220_73640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8585 n_85500_82040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8586 n_68780_82040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8587 n_71060_82040 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8588 n_60040_56840 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8589 n_60040_59640 0 PWL(70000ps 0uA 70030ps 0uA 70031ps 30uA 70059ps 30uA 70060ps 0uA)
I8590 n_91960_87640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8591 n_87020_87640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8592 n_93100_87640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8593 n_90440_62440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8594 n_83600_87640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8595 n_84740_87640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8596 n_54720_48440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8597 n_44080_54040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8598 n_40660_56840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8599 n_79040_42840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8600 n_48640_40040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8601 n_50920_48440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8602 n_63840_40040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8603 n_91580_40040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8604 n_56620_40040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8605 n_67260_40040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8606 n_46360_40040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8607 n_40280_40040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8608 n_60040_45640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8609 n_72200_40040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8610 n_82080_48440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8611 n_77140_40040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8612 n_55100_40040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8613 n_43320_59640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8614 n_42180_73640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8615 n_44460_68040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8616 n_46740_65240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8617 n_52060_73640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8618 n_46740_59640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8619 n_54720_42840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8620 n_74860_40040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8621 n_80180_45640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8622 n_71820_42840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8623 n_56620_45640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8624 n_41420_40040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8625 n_49400_40040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8626 n_66880_45640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8627 n_57760_40040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8628 n_92720_40040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8629 n_63460_42840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8630 n_51680_48440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8631 n_47880_42840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8632 n_78280_48440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8633 n_41420_54040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8634 n_49020_51240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8635 n_54720_51240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8636 n_81700_87640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8637 n_80180_87640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8638 n_90820_59640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8639 n_90060_87640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8640 n_85120_84840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8641 n_87400_84840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8642 n_68780_79240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8643 n_88920_82040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8644 n_82080_84840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8645 n_85880_87640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8646 n_89300_59640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8647 n_80560_84840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8648 n_81700_82040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8649 n_80180_59640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8650 n_82080_56840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8651 n_78660_56840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8652 n_76760_65240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8653 n_80940_62440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8654 n_76760_56840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8655 n_78660_65240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8656 n_77900_68040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8657 n_79040_68040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8658 n_78280_70840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8659 n_73720_73640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8660 n_70300_79240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8661 n_71820_79240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8662 n_88920_79240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8663 n_70300_84840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8664 n_73720_82040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8665 n_85500_56840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8666 n_82080_59640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8667 n_83600_59640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8668 n_76760_79240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8669 n_80560_79240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8670 n_74860_84840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8671 n_76760_82040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8672 n_70300_51240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8673 n_50920_51240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8674 n_52060_51240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8675 n_79040_51240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8676 n_51680_45640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8677 n_53200_48440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8678 n_65360_42840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8679 n_92720_42840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8680 n_61560_40040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8681 n_68020_48440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8682 n_51300_40040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8683 n_43320_40040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8684 n_53200_45640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8685 n_73720_45640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8686 n_82080_45640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8687 n_73340_40040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8688 n_53200_42840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8689 n_58900_48440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8690 n_57000_54040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8691 n_49780_56840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8692 n_48260_62440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8693 n_52060_54040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8694 n_48260_65240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8695 n_49780_62440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8696 n_44840_73640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8697 n_50920_68040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8698 n_72200_56840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8699 n_56620_65240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8700 n_58520_65240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8701 n_60420_65240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8702 n_73720_62440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8703 n_76380_62440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8704 n_63080_82040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8705 n_75240_59640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8706 n_77520_62440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8707 n_73340_59640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8708 n_55100_70840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8709 n_53580_70840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8710 n_50920_70840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8711 n_50920_73640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8712 n_46740_73640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8713 n_46360_76440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8714 n_48260_73640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8715 n_61560_73640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8716 n_66880_73640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8717 n_63460_70840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8718 n_74100_68040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8719 n_65360_70840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8720 n_68780_68040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8721 n_75240_65240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8722 n_68020_62440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8723 n_68780_70840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8724 n_53580_65240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8725 n_53580_68040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8726 n_49400_70840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8727 n_46740_70840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8728 n_48260_76440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8729 n_58520_70840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8730 n_60420_70840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8731 n_63080_73640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8732 n_71820_73640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8733 n_76760_73640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8734 n_67260_70840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8735 n_58140_51240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8736 n_65740_73640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8737 n_70300_76440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8738 n_47500_56840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8739 n_52820_79240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8740 n_61940_84840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8741 n_63080_84840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8742 n_52440_87640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8743 n_49400_87640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8744 n_64220_82040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8745 n_58140_87640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8746 n_46740_51240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8747 n_66880_62440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8748 n_65360_54040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8749 n_63080_54040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8750 n_54340_87640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8751 n_67260_82040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8752 n_53580_87640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8753 n_58520_84840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8754 n_64600_84840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8755 n_73340_87640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8756 n_63460_87640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8757 n_67260_65240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8758 n_63460_62440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8759 n_60040_54040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8760 n_66880_59640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8761 n_70300_59640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8762 n_70300_56840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8763 n_71820_59640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8764 n_71820_70840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8765 n_55100_79240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8766 n_59660_82040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8767 n_56240_82040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8768 n_87400_62440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8769 n_87020_59640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8770 n_84740_68040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8771 n_85880_73640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8772 n_83600_76440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8773 n_85500_76440 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8774 n_85500_79240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8775 n_87400_82040 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8776 n_83600_79240 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8777 n_44460_56840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8778 n_60040_56840 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8779 n_60040_59640 0 PWL(72000ps 0uA 72030ps 0uA 72031ps 30uA 72059ps 30uA 72060ps 0uA)
I8780 n_90820_68040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8781 n_91200_70840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8782 n_87020_87640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8783 n_93480_76440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8784 n_93100_84840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8785 n_65740_40040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8786 n_40280_54040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8787 n_44080_54040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8788 n_63840_45640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8789 n_79040_42840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8790 n_48640_40040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8791 n_70300_40040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8792 n_91580_40040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8793 n_52440_40040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8794 n_90440_40040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8795 n_93480_45640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8796 n_80560_40040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8797 n_40280_40040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8798 n_40280_48440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8799 n_72200_40040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8800 n_79040_40040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8801 n_82080_48440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8802 n_77140_40040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8803 n_40660_45640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8804 n_40660_51240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8805 n_43320_59640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8806 n_50160_59640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8807 n_42180_73640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8808 n_45600_68040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8809 n_43320_62440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8810 n_40660_65240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8811 n_41800_68040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8812 n_44460_62440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8813 n_47500_68040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8814 n_52060_73640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8815 n_51300_59640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8816 n_46740_59640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8817 n_44840_51240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8818 n_45220_48440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8819 n_74860_40040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8820 n_80180_45640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8821 n_76760_42840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8822 n_71820_42840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8823 n_41420_48440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8824 n_41420_40040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8825 n_80180_42840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8826 n_88920_45640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8827 n_83600_42840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8828 n_51680_42840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8829 n_92720_40040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8830 n_68400_40040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8831 n_47880_42840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8832 n_78280_48440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8833 n_64980_48440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8834 n_49020_51240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8835 n_47880_54040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8836 n_63080_51240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8837 n_90820_84840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8838 n_90440_76440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8839 n_85120_84840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8840 n_87400_73640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8841 n_88540_68040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8842 n_87400_65240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8843 n_87400_76440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8844 n_82080_84840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8845 n_87400_56840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8846 n_90820_56840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8847 n_77520_54040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8848 n_87400_79240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8849 n_89300_59640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8850 n_92720_59640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8851 n_88920_65240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8852 n_91960_68040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8853 n_88920_76440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8854 n_90820_82040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8855 n_81700_82040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8856 n_79040_87640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8857 n_79040_54040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8858 n_80560_54040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8859 n_80560_56840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8860 n_80180_59640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8861 n_78660_56840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8862 n_83600_56840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8863 n_76380_54040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8864 n_76760_65240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8865 n_80940_62440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8866 n_76760_56840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8867 n_78660_65240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8868 n_80560_65240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8869 n_76000_70840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8870 n_79040_68040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8871 n_78280_70840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8872 n_75240_73640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8873 n_73720_79240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8874 n_70300_79240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8875 n_71820_79240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8876 n_88920_79240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8877 n_70300_84840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8878 n_73720_82040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8879 n_85500_56840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8880 n_86260_54040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8881 n_82080_59640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8882 n_85500_59640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8883 n_84740_65240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8884 n_83600_59640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8885 n_85880_65240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8886 n_87400_68040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8887 n_80560_70840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8888 n_80560_73640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8889 n_76760_82040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8890 n_67260_51240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8891 n_71820_51240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8892 n_71820_54040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8893 n_53200_51240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8894 n_70300_51240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8895 n_53580_54040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8896 n_68020_54040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8897 n_59280_51240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8898 n_61940_51240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8899 n_46360_54040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8900 n_47880_51240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8901 n_41800_56840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8902 n_52060_51240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8903 n_70300_54040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8904 n_61560_54040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8905 n_66120_51240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8906 n_79040_51240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8907 n_51680_45640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8908 n_70300_42840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8909 n_92720_42840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8910 n_50540_42840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8911 n_85500_42840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8912 n_88920_42840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8913 n_82080_42840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8914 n_43320_40040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8915 n_42940_48440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8916 n_73720_45640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8917 n_76760_45640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8918 n_82080_45640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8919 n_73340_40040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8920 n_44080_48440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8921 n_43320_51240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8922 n_57000_54040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8923 n_61940_59640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8924 n_49780_56840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8925 n_51680_56840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8926 n_48260_65240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8927 n_59660_62440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8928 n_50920_68040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8929 n_53580_59640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8930 n_53580_56840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8931 n_49400_65240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8932 n_56620_65240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8933 n_58520_65240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8934 n_60420_65240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8935 n_73720_62440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8936 n_75240_62440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8937 n_76380_59640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8938 n_55100_56840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8939 n_55100_70840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8940 n_53580_70840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8941 n_50920_70840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8942 n_46360_76440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8943 n_40660_76440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8944 n_48260_73640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8945 n_40660_70840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8946 n_61560_73640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8947 n_66880_73640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8948 n_55480_48440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8949 n_68780_70840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8950 n_56240_59640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8951 n_53580_68040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8952 n_49400_70840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8953 n_48260_76440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8954 n_58520_70840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8955 n_60420_70840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8956 n_63080_73640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8957 n_67260_70840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8958 n_46360_68040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8959 n_48260_56840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8960 n_41800_70840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8961 n_40280_82040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8962 n_40280_87640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8963 n_50920_82040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8964 n_53580_82040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8965 n_52820_79240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8966 n_44080_59640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8967 n_42940_56840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8968 n_40280_84840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8969 n_41420_87640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8970 n_46740_87640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8971 n_46740_84840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8972 n_49400_84840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8973 n_52440_87640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8974 n_49400_87640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8975 n_64220_82040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8976 n_58140_87640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8977 n_55100_82040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8978 n_42940_54040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8979 n_46740_51240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8980 n_43320_68040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8981 n_44080_65240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8982 n_65360_62440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8983 n_65360_54040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8984 n_65360_56840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8985 n_63080_54040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8986 n_54340_87640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8987 n_67260_82040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8988 n_53580_87640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8989 n_57000_87640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8990 n_60040_54040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8991 n_70300_59640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8992 n_70300_56840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8993 n_71820_59640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8994 n_71820_70840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8995 n_55100_79240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8996 n_59660_82040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8997 n_56240_82040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8998 n_88160_59640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I8999 n_85880_62440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I9000 n_83220_65240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I9001 n_84740_62440 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I9002 n_83220_68040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I9003 n_84740_68040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I9004 n_83600_70840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I9005 n_85500_70840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I9006 n_84740_73640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I9007 n_85880_68040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I9008 n_85880_73640 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I9009 n_83600_82040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I9010 n_83600_79240 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I9011 n_69920_82040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I9012 n_71060_82040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I9013 n_72200_82040 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I9014 n_61560_56840 0 PWL(74000ps 0uA 74030ps 0uA 74031ps 30uA 74059ps 30uA 74060ps 0uA)
I9015 n_93480_62440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9016 n_91200_70840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9017 n_93480_79240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9018 n_91960_87640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9019 n_93480_56840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9020 n_90440_62440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9021 n_93100_84840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9022 n_83600_87640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9023 n_84740_87640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9024 n_54720_48440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9025 n_61940_48440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9026 n_40280_54040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9027 n_40660_56840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9028 n_92340_48440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9029 n_50920_48440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9030 n_70300_40040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9031 n_87020_40040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9032 n_52440_40040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9033 n_56620_40040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9034 n_90440_40040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9035 n_93480_45640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9036 n_46360_40040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9037 n_40280_48440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9038 n_72200_40040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9039 n_79040_40040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9040 n_40660_51240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9041 n_43320_59640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9042 n_42180_73640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9043 n_45600_68040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9044 n_43320_62440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9045 n_44460_62440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9046 n_47500_68040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9047 n_52060_73640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9048 n_46740_59640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9049 n_44840_51240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9050 n_76760_42840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9051 n_71820_42840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9052 n_41420_48440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9053 n_49400_40040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9054 n_88920_45640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9055 n_83600_42840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9056 n_57760_40040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9057 n_51680_42840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9058 n_87020_45640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9059 n_68400_40040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9060 n_51680_48440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9061 n_85120_48440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9062 n_41420_54040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9063 n_47880_54040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9064 n_60040_48440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9065 n_54720_51240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9066 n_81700_87640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9067 n_80180_87640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9068 n_90820_84840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9069 n_90820_59640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9070 n_88920_56840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9071 n_87400_84840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9072 n_91580_79240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9073 n_87400_73640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9074 n_91580_62440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9075 n_90820_65240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9076 n_87400_76440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9077 n_92340_76440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9078 n_88920_82040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9079 n_90820_56840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9080 n_77520_54040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9081 n_87400_79240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9082 n_92720_59640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9083 n_88920_65240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9084 n_91960_68040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9085 n_90820_82040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9086 n_80560_84840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9087 n_79040_87640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9088 n_79040_54040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9089 n_80560_54040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9090 n_80560_56840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9091 n_82080_56840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9092 n_83600_56840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9093 n_80560_65240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9094 n_77900_68040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9095 n_76000_70840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9096 n_75240_73640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9097 n_75240_76440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9098 n_73720_79240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9099 n_73720_73640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9100 n_70300_79240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9101 n_71820_79240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9102 n_88920_79240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9103 n_82080_59640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9104 n_82080_65240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9105 n_80560_70840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9106 n_80560_73640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9107 n_72200_76440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9108 n_76760_79240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9109 n_80560_79240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9110 n_71820_51240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9111 n_71820_54040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9112 n_53200_51240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9113 n_53580_54040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9114 n_68020_54040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9115 n_59280_51240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9116 n_46360_54040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9117 n_47880_51240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9118 n_50920_51240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9119 n_41800_56840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9120 n_70300_54040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9121 n_61560_54040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9122 n_83600_48440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9123 n_53200_48440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9124 n_70300_42840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9125 n_90440_45640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9126 n_50540_42840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9127 n_61560_40040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9128 n_85500_42840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9129 n_88920_42840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9130 n_51300_40040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9131 n_42940_48440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9132 n_73720_45640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9133 n_76760_45640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9134 n_43320_51240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9135 n_61940_59640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9136 n_49780_56840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9137 n_51680_56840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9138 n_52060_54040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9139 n_59660_62440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9140 n_53580_56840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9141 n_53580_62440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9142 n_52060_65240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9143 n_77520_62440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9144 n_55100_70840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9145 n_53580_70840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9146 n_50920_70840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9147 n_66880_73640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9148 n_58140_79240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9149 n_55480_48440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9150 n_68780_70840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9151 n_56240_59640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9152 n_53580_68040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9153 n_49400_70840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9154 n_48640_79240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9155 n_60040_76440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9156 n_56620_79240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9157 n_63080_79240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9158 n_61560_79240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9159 n_52060_82040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9160 n_65740_76440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9161 n_67260_70840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9162 n_58140_51240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9163 n_70300_48440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9164 n_46360_68040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9165 n_48260_56840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9166 n_41800_70840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9167 n_40660_79240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9168 n_43700_79240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9169 n_44080_84840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9170 n_63080_76440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9171 n_80560_76440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9172 n_50920_82040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9173 n_49400_82040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9174 n_47120_82040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9175 n_53580_82040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9176 n_50160_84840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9177 n_65740_73640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9178 n_47500_56840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9179 n_52820_79240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9180 n_44080_59640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9181 n_42940_56840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9182 n_40280_84840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9183 n_49400_84840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9184 n_52440_87640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9185 n_58140_87640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9186 n_55100_82040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9187 n_46740_51240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9188 n_44080_65240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9189 n_43320_76440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9190 n_41800_82040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9191 n_65360_62440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9192 n_65360_54040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9193 n_65360_56840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9194 n_63080_54040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9195 n_45220_87640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9196 n_51680_84840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9197 n_54340_87640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9198 n_53580_87640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9199 n_73340_87640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9200 n_57000_87640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9201 n_60040_54040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9202 n_71820_70840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9203 n_67260_76440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9204 n_65740_79240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9205 n_64600_79240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9206 n_57380_82040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9207 n_55100_79240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9208 n_58520_82040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9209 n_56240_82040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9210 n_88160_59640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9211 n_85880_62440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9212 n_83220_65240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9213 n_84740_62440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9214 n_84740_73640 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9215 n_83600_76440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9216 n_85500_76440 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9217 n_85500_79240 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9218 n_87400_82040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9219 n_83600_82040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9220 n_69920_82040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9221 n_71060_82040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9222 n_72200_82040 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9223 n_61560_56840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9224 n_44460_56840 0 PWL(76000ps 0uA 76030ps 0uA 76031ps 30uA 76059ps 30uA 76060ps 0uA)
I9225 n_92340_54040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9226 n_91200_70840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9227 n_93480_79240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9228 n_87020_87640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9229 n_93100_87640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9230 n_93480_56840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9231 n_93480_73640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9232 n_84740_87640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9233 n_65740_40040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9234 n_65740_45640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9235 n_40660_56840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9236 n_63840_45640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9237 n_93480_54040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9238 n_50920_48440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9239 n_63840_40040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9240 n_70300_40040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9241 n_91580_40040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9242 n_87020_40040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9243 n_52440_40040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9244 n_40660_42840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9245 n_56620_40040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9246 n_67260_40040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9247 n_80560_40040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9248 n_40280_48440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9249 n_60040_45640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9250 n_82080_48440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9251 n_77140_40040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9252 n_55100_40040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9253 n_40660_45640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9254 n_50160_59640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9255 n_42180_73640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9256 n_44460_68040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9257 n_46740_65240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9258 n_52060_73640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9259 n_51300_59640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9260 n_45220_48440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9261 n_54720_42840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9262 n_74860_40040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9263 n_80180_45640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9264 n_56620_45640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9265 n_41420_48440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9266 n_80180_42840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9267 n_66880_45640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9268 n_57760_40040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9269 n_43700_42840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9270 n_51680_42840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9271 n_87020_45640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9272 n_92720_40040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9273 n_68400_40040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9274 n_63460_42840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9275 n_51680_48440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9276 n_92340_51240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9277 n_64980_48440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9278 n_41420_54040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9279 n_64600_51240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9280 n_63080_51240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9281 n_81700_87640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9282 n_90440_73640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9283 n_88920_56840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9284 n_90060_87640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9285 n_85120_84840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9286 n_91580_79240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9287 n_87400_73640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9288 n_89300_54040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9289 n_88920_51240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9290 n_87400_76440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9291 n_92340_76440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9292 n_82080_84840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9293 n_85880_87640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9294 n_87400_56840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9295 n_89300_73640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9296 n_81700_82040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9297 n_80180_59640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9298 n_76380_54040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9299 n_80560_65240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9300 n_77900_68040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9301 n_76000_70840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9302 n_79040_68040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9303 n_78280_70840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9304 n_75240_73640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9305 n_74860_70840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9306 n_73720_70840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9307 n_75240_76440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9308 n_73720_79240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9309 n_73720_73640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9310 n_70300_79240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9311 n_67260_84840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9312 n_88920_79240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9313 n_67260_87640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9314 n_68780_87640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9315 n_68780_84840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9316 n_70300_84840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9317 n_72200_84840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9318 n_87400_48440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9319 n_80560_73640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9320 n_78660_79240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9321 n_76760_76440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9322 n_78280_82040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9323 n_80180_82040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9324 n_76760_84840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9325 n_76380_87640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9326 n_74860_84840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9327 n_76760_82040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9328 n_67260_51240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9329 n_68780_51240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9330 n_52060_51240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9331 n_66120_51240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9332 n_90820_51240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9333 n_53200_48440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9334 n_65360_42840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9335 n_70300_42840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9336 n_92720_42840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9337 n_90440_45640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9338 n_50540_42840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9339 n_45220_42840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9340 n_61560_40040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9341 n_68020_48440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9342 n_82080_42840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9343 n_42940_48440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9344 n_53200_45640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9345 n_82080_45640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9346 n_73340_40040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9347 n_53200_42840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9348 n_44080_48440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9349 n_58900_48440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9350 n_57000_54040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9351 n_52060_54040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9352 n_48260_65240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9353 n_59660_62440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9354 n_50920_68040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9355 n_53580_59640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9356 n_53580_62440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9357 n_52060_65240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9358 n_49400_65240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9359 n_56620_65240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9360 n_61560_62440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9361 n_61560_65240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9362 n_59660_68040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9363 n_60800_68040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9364 n_60040_73640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9365 n_63080_65240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9366 n_61940_68040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9367 n_59660_70840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9368 n_55100_56840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9369 n_55100_70840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9370 n_53580_70840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9371 n_50920_70840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9372 n_50920_73640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9373 n_49400_73640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9374 n_55860_68040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9375 n_46360_76440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9376 n_48260_73640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9377 n_49780_76440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9378 n_50920_79240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9379 n_58520_73640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9380 n_70300_73640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9381 n_55480_48440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9382 n_53580_65240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9383 n_53580_68040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9384 n_49400_70840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9385 n_46740_70840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9386 n_48260_76440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9387 n_47500_79240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9388 n_58520_70840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9389 n_60420_70840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9390 n_71820_73640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9391 n_80560_76440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9392 n_47500_56840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9393 n_50920_87640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9394 n_59660_84840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9395 n_42940_54040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9396 n_44080_82040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9397 n_41800_82040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9398 n_65360_62440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9399 n_65360_54040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9400 n_65360_56840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9401 n_68780_56840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9402 n_59280_87640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9403 n_51680_84840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9404 n_74860_87640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9405 n_54340_87640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9406 n_58520_84840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9407 n_56240_76440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9408 n_65360_65240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9409 n_63460_62440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9410 n_63460_59640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9411 n_63460_56840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9412 n_67260_56840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9413 n_70300_59640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9414 n_70300_56840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9415 n_71820_59640 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9416 n_70300_65240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9417 n_71820_65240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9418 n_71820_68040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9419 n_70300_70840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9420 n_71820_70840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9421 n_56620_84840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9422 n_87400_62440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9423 n_88920_62440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9424 n_83220_62440 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9425 n_83220_68040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9426 n_83600_70840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9427 n_85500_70840 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9428 n_85880_68040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9429 n_85500_82040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9430 n_68780_82040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9431 n_71060_82040 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9432 n_43320_65240 0 PWL(78000ps 0uA 78030ps 0uA 78031ps 30uA 78059ps 30uA 78060ps 0uA)
I9433 n_90820_68040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9434 n_93480_79240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9435 n_91960_87640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9436 n_90440_62440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9437 n_93480_68040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9438 n_93480_73640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9439 n_83600_87640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9440 n_84740_87640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9441 n_56240_48440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9442 n_40280_54040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9443 n_44080_54040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9444 n_40660_56840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9445 n_93480_48440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9446 n_41800_42840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9447 n_48640_40040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9448 n_50920_48440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9449 n_63840_40040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9450 n_40660_42840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9451 n_67260_40040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9452 n_93480_45640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9453 n_80560_40040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9454 n_40280_48440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9455 n_79040_40040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9456 n_55100_40040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9457 n_40660_51240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9458 n_50160_59640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9459 n_42180_73640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9460 n_40660_65240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9461 n_41800_68040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9462 n_52060_73640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9463 n_51300_59640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9464 n_44840_51240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9465 n_54720_42840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9466 n_76760_42840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9467 n_41420_48440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9468 n_80180_42840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9469 n_88920_45640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9470 n_66880_45640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9471 n_43700_42840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9472 n_63460_42840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9473 n_51680_48440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9474 n_47880_42840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9475 n_48260_45640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9476 n_90440_48440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9477 n_41420_54040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9478 n_49020_51240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9479 n_47880_54040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9480 n_55100_54040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9481 n_81700_87640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9482 n_80180_87640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9483 n_90440_73640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9484 n_92340_65240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9485 n_90820_59640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9486 n_87400_84840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9487 n_91580_79240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9488 n_88540_68040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9489 n_87780_54040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9490 n_88920_51240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9491 n_83220_54040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9492 n_91200_54040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9493 n_87400_65240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9494 n_87400_70840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9495 n_87400_76440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9496 n_92340_76440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9497 n_87780_87640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9498 n_83600_51240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9499 n_80560_51240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9500 n_84740_54040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9501 n_87400_56840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9502 n_90820_56840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9503 n_77520_54040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9504 n_87400_79240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9505 n_92720_59640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9506 n_88920_65240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9507 n_89300_73640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9508 n_80560_84840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9509 n_81700_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9510 n_79040_54040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9511 n_80560_54040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9512 n_82080_54040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9513 n_80180_59640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9514 n_79040_68040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9515 n_65740_84840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9516 n_62320_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9517 n_70300_87640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9518 n_73720_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9519 n_72200_84840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9520 n_85500_56840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9521 n_85500_59640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9522 n_84740_65240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9523 n_82080_68040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9524 n_87400_68040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9525 n_82080_70840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9526 n_77140_70840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9527 n_81700_73640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9528 n_80560_73640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9529 n_78660_73640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9530 n_79040_70840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9531 n_78660_79240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9532 n_76760_76440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9533 n_78280_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9534 n_80560_79240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9535 n_80180_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9536 n_76760_84840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9537 n_76380_87640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9538 n_74860_84840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9539 n_74860_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9540 n_76760_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9541 n_68020_54040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9542 n_49780_54040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9543 n_50920_51240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9544 n_52060_51240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9545 n_87400_51240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9546 n_49400_48440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9547 n_51680_45640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9548 n_53200_48440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9549 n_65360_42840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9550 n_45220_42840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9551 n_68020_48440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9552 n_88920_42840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9553 n_82080_42840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9554 n_42940_48440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9555 n_76760_45640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9556 n_53200_42840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9557 n_43320_51240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9558 n_57000_54040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9559 n_48260_65240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9560 n_59660_62440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9561 n_50920_68040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9562 n_53580_59640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9563 n_53580_62440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9564 n_52060_65240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9565 n_49400_65240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9566 n_56620_65240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9567 n_61560_62440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9568 n_61560_65240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9569 n_59660_68040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9570 n_60800_68040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9571 n_63460_68040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9572 n_60040_73640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9573 n_63080_65240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9574 n_61940_68040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9575 n_59660_70840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9576 n_55100_70840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9577 n_53580_70840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9578 n_50920_70840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9579 n_50920_73640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9580 n_49400_73640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9581 n_46740_73640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9582 n_46360_76440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9583 n_40660_76440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9584 n_40660_70840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9585 n_58520_68040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9586 n_61560_73640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9587 n_58140_79240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9588 n_74100_68040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9589 n_75240_65240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9590 n_55480_48440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9591 n_48260_76440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9592 n_47500_79240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9593 n_48640_79240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9594 n_58520_70840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9595 n_60040_76440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9596 n_60420_70840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9597 n_63080_73640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9598 n_60040_79240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9599 n_61560_79240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9600 n_52060_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9601 n_58140_51240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9602 n_40660_79240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9603 n_40280_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9604 n_43700_79240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9605 n_44080_84840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9606 n_40280_87640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9607 n_57380_76440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9608 n_80560_76440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9609 n_50920_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9610 n_54720_84840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9611 n_47120_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9612 n_53580_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9613 n_50160_84840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9614 n_52820_79240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9615 n_41420_87640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9616 n_46740_87640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9617 n_61940_84840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9618 n_49400_84840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9619 n_49400_87640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9620 n_64220_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9621 n_50920_87640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9622 n_59660_84840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9623 n_55100_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9624 n_43320_68040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9625 n_43320_76440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9626 n_44080_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9627 n_65360_62440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9628 n_65360_54040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9629 n_65360_56840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9630 n_68780_56840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9631 n_45220_87640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9632 n_59280_87640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9633 n_74860_87640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9634 n_54340_87640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9635 n_67260_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9636 n_58520_84840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9637 n_56240_76440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9638 n_65360_65240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9639 n_63460_62440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9640 n_63460_59640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9641 n_63460_56840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9642 n_67260_56840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9643 n_66880_59640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9644 n_70300_59640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9645 n_70300_56840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9646 n_71820_59640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9647 n_70300_65240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9648 n_68400_65240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9649 n_71820_65240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9650 n_71820_68040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9651 n_70300_70840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9652 n_67260_76440 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9653 n_65740_79240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9654 n_64600_79240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9655 n_57380_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9656 n_58520_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9657 n_59660_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9658 n_56620_84840 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9659 n_87020_59640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9660 n_84740_68040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9661 n_85880_73640 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9662 n_81700_79240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9663 n_85500_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9664 n_68780_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9665 n_71060_82040 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9666 n_43320_65240 0 PWL(80000ps 0uA 80030ps 0uA 80031ps 30uA 80059ps 30uA 80060ps 0uA)
I9667 n_93480_62440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9668 n_93480_79240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9669 n_90440_62440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9670 n_93480_73640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9671 n_40280_54040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9672 n_41800_42840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9673 n_70300_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9674 n_91580_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9675 n_87020_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9676 n_88160_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9677 n_56620_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9678 n_67260_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9679 n_90440_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9680 n_93480_45640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9681 n_80560_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9682 n_46360_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9683 n_40280_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9684 n_60040_45640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9685 n_72200_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9686 n_55100_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9687 n_40660_45640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9688 n_40660_51240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9689 n_50160_59640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9690 n_51300_59640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9691 n_44840_51240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9692 n_45220_48440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9693 n_54720_42840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9694 n_71820_42840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9695 n_56620_45640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9696 n_41420_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9697 n_49400_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9698 n_80180_42840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9699 n_88920_45640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9700 n_83600_42840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9701 n_66880_45640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9702 n_57760_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9703 n_83600_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9704 n_87020_45640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9705 n_92720_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9706 n_68400_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9707 n_48260_45640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9708 n_47880_54040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9709 n_90440_73640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9710 n_90820_59640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9711 n_91580_79240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9712 n_91580_62440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9713 n_87780_54040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9714 n_88920_51240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9715 n_83220_54040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9716 n_91200_54040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9717 n_90820_65240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9718 n_87400_70840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9719 n_87400_76440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9720 n_92340_76440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9721 n_87780_87640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9722 n_88920_82040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9723 n_83600_51240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9724 n_80560_51240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9725 n_84740_54040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9726 n_87400_56840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9727 n_90820_56840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9728 n_77520_54040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9729 n_87400_79240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9730 n_92720_59640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9731 n_89300_73640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9732 n_79040_54040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9733 n_80560_54040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9734 n_82080_54040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9735 n_80560_65240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9736 n_77900_68040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9737 n_76000_70840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9738 n_75240_73640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9739 n_74860_70840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9740 n_73720_79240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9741 n_70300_79240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9742 n_67260_84840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9743 n_67260_87640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9744 n_65740_84840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9745 n_62320_82040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9746 n_68780_87640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9747 n_71820_87640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9748 n_85500_56840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9749 n_82080_59640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9750 n_85500_59640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9751 n_84740_65240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9752 n_82080_65240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9753 n_82080_68040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9754 n_82080_70840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9755 n_81700_73640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9756 n_80560_73640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9757 n_78660_73640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9758 n_79040_70840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9759 n_76760_76440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9760 n_76760_79240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9761 n_74860_84840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9762 n_74860_82040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9763 n_76760_82040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9764 n_49780_54040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9765 n_49400_48440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9766 n_70300_42840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9767 n_92720_42840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9768 n_90440_45640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9769 n_85500_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9770 n_61560_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9771 n_68020_48440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9772 n_85500_42840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9773 n_88920_42840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9774 n_82080_42840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9775 n_51300_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9776 n_43320_40040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9777 n_53200_45640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9778 n_73720_45640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9779 n_53200_42840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9780 n_44080_48440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9781 n_43320_51240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9782 n_58900_48440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9783 n_57000_54040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9784 n_48260_65240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9785 n_50920_68040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9786 n_72200_56840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9787 n_53580_59640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9788 n_53580_62440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9789 n_52060_65240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9790 n_49400_65240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9791 n_56620_65240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9792 n_58520_65240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9793 n_60420_65240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9794 n_73720_62440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9795 n_60040_73640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9796 n_75240_62440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9797 n_76380_59640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9798 n_75240_59640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9799 n_72200_62440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9800 n_61940_68040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9801 n_59660_70840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9802 n_55860_68040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9803 n_46360_79240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9804 n_61560_73640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9805 n_66880_73640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9806 n_55480_48440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9807 n_68780_70840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9808 n_48260_76440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9809 n_47500_79240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9810 n_45600_84840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9811 n_48640_79240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9812 n_58520_70840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9813 n_49400_79240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9814 n_60040_76440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9815 n_60420_70840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9816 n_63080_73640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9817 n_56620_79240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9818 n_65740_76440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9819 n_67260_70840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9820 n_58140_51240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9821 n_70300_48440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9822 n_57380_76440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9823 n_80560_76440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9824 n_49400_82040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9825 n_54720_84840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9826 n_65740_73640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9827 n_47500_56840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9828 n_41420_87640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9829 n_46740_87640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9830 n_43320_87640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9831 n_61940_84840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9832 n_52440_87640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9833 n_58140_87640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9834 n_42940_54040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9835 n_46740_51240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9836 n_45220_87640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9837 n_59280_87640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9838 n_51680_84840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9839 n_60800_84840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9840 n_61180_82040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9841 n_54340_76440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9842 n_54340_87640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9843 n_53580_87640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9844 n_57000_87640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9845 n_71820_65240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9846 n_73720_65240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9847 n_68780_76440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9848 n_55100_79240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9849 n_56240_82040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9850 n_83220_62440 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9851 n_83600_70840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9852 n_83220_73640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9853 n_85880_73640 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9854 n_81700_79240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9855 n_68780_82040 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9856 n_43320_65240 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9857 n_44460_56840 0 PWL(82000ps 0uA 82030ps 0uA 82031ps 30uA 82059ps 30uA 82060ps 0uA)
I9858 n_90820_68040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9859 n_91200_70840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9860 n_93480_79240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9861 n_91960_87640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9862 n_87020_87640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9863 n_93480_68040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9864 n_93480_73640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9865 n_93480_76440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9866 n_93100_84840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9867 n_84740_87640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9868 n_54720_48440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9869 n_56240_48440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9870 n_65740_45640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9871 n_44080_54040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9872 n_79040_42840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9873 n_93480_48440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9874 n_93480_54040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9875 n_48640_40040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9876 n_91580_40040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9877 n_42940_42840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9878 n_56620_40040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9879 n_80560_40040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9880 n_72200_40040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9881 n_40660_45640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9882 n_40660_51240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9883 n_44460_68040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9884 n_45600_68040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9885 n_43320_62440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9886 n_44460_62440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9887 n_47500_68040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9888 n_46740_65240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9889 n_44840_51240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9890 n_45220_48440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9891 n_71820_42840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9892 n_80180_42840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9893 n_57760_40040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9894 n_44840_45640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9895 n_92720_40040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9896 n_47880_42840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9897 n_92340_51240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9898 n_90440_48440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9899 n_78280_48440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9900 n_49020_51240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9901 n_64600_51240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9902 n_55100_54040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9903 n_54720_51240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9904 n_81700_87640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9905 n_90820_84840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9906 n_90440_76440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9907 n_90440_73640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9908 n_92340_65240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9909 n_85120_84840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9910 n_87400_84840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9911 n_91580_79240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9912 n_87400_73640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9913 n_88540_68040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9914 n_68780_79240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9915 n_87780_54040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9916 n_88920_51240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9917 n_83220_54040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9918 n_91200_54040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9919 n_92340_56840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9920 n_90820_65240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9921 n_88920_70840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9922 n_87400_76440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9923 n_92340_76440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9924 n_88920_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9925 n_83600_84840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9926 n_83600_51240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9927 n_80560_51240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9928 n_84740_54040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9929 n_87400_56840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9930 n_90820_56840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9931 n_77520_54040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9932 n_87400_79240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9933 n_91960_68040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9934 n_89300_73640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9935 n_90060_79240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9936 n_90820_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9937 n_79040_87640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9938 n_79040_54040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9939 n_80560_54040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9940 n_82080_54040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9941 n_80560_56840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9942 n_82080_56840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9943 n_78660_56840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9944 n_80940_62440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9945 n_76760_56840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9946 n_78280_70840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9947 n_73720_70840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9948 n_75240_76440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9949 n_88920_79240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9950 n_68780_84840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9951 n_71820_87640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9952 n_70300_87640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9953 n_70300_84840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9954 n_73720_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9955 n_85500_56840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9956 n_82080_59640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9957 n_85500_59640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9958 n_84740_65240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9959 n_83600_59640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9960 n_82080_65240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9961 n_85880_65240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9962 n_77140_70840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9963 n_80560_73640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9964 n_74860_84840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9965 n_76760_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9966 n_70300_51240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9967 n_68020_54040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9968 n_68780_51240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9969 n_50920_51240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9970 n_79040_51240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9971 n_87400_51240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9972 n_90820_51240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9973 n_51680_45640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9974 n_92720_42840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9975 n_46740_45640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9976 n_61560_40040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9977 n_82080_42840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9978 n_73720_45640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9979 n_44080_48440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9980 n_43320_51240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9981 n_57000_54040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9982 n_63460_68040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9983 n_60040_73640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9984 n_76380_59640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9985 n_63080_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9986 n_77520_62440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9987 n_72200_62440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9988 n_73340_59640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9989 n_61940_68040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9990 n_59660_70840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9991 n_46740_73640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9992 n_40660_76440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9993 n_48260_73640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9994 n_40660_70840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9995 n_49780_76440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9996 n_50920_79240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9997 n_46360_79240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9998 n_58520_68040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I9999 n_58520_73640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10000 n_70300_73640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10001 n_66880_73640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10002 n_58140_79240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10003 n_63460_70840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10004 n_65360_70840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10005 n_68780_68040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10006 n_68020_62440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10007 n_55480_48440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10008 n_68780_70840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10009 n_53580_65240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10010 n_53580_68040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10011 n_49400_70840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10012 n_46740_70840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10013 n_48260_76440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10014 n_47500_79240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10015 n_45600_84840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10016 n_48640_79240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10017 n_58520_70840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10018 n_49400_79240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10019 n_60040_76440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10020 n_60420_70840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10021 n_76760_73640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10022 n_56620_79240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10023 n_60040_79240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10024 n_63080_79240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10025 n_61560_79240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10026 n_52060_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10027 n_65740_76440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10028 n_68400_73640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10029 n_58140_51240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10030 n_70300_48440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10031 n_46360_68040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10032 n_44840_70840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10033 n_43320_70840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10034 n_41800_70840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10035 n_40280_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10036 n_40280_87640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10037 n_63080_76440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10038 n_50920_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10039 n_49400_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10040 n_54720_84840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10041 n_47120_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10042 n_53580_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10043 n_50160_84840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10044 n_65740_73640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10045 n_47500_56840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10046 n_44080_59640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10047 n_42940_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10048 n_42940_84840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10049 n_40280_84840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10050 n_46740_87640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10051 n_61940_84840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10052 n_49400_84840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10053 n_52440_87640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10054 n_49400_87640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10055 n_64220_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10056 n_59660_84840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10057 n_55100_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10058 n_42940_54040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10059 n_46740_51240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10060 n_66880_62440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10061 n_65360_54040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10062 n_63080_54040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10063 n_60800_84840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10064 n_61180_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10065 n_54340_87640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10066 n_67260_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10067 n_58520_84840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10068 n_73340_87640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10069 n_57000_87640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10070 n_63460_87640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10071 n_67260_65240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10072 n_63460_62440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10073 n_60040_54040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10074 n_71820_59640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10075 n_68400_65240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10076 n_71820_65240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10077 n_73720_65240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10078 n_71820_70840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10079 n_68780_76440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10080 n_58520_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10081 n_59660_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10082 n_56240_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10083 n_83220_62440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10084 n_84740_68040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10085 n_83600_70840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10086 n_83220_73640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10087 n_85880_73640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10088 n_83600_76440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10089 n_85500_76440 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10090 n_85500_79240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10091 n_87400_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10092 n_83600_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10093 n_83600_79240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10094 n_69920_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10095 n_68780_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10096 n_71060_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10097 n_72200_82040 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10098 n_43320_65240 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10099 n_60040_56840 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10100 n_60040_59640 0 PWL(84000ps 0uA 84030ps 0uA 84031ps 30uA 84059ps 30uA 84060ps 0uA)
I10101 n_92340_54040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10102 n_90820_68040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10103 n_91200_70840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10104 n_93480_79240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10105 n_90440_62440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10106 n_93480_76440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10107 n_65740_40040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10108 n_54720_48440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10109 n_65740_45640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10110 n_63840_45640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10111 n_79040_42840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10112 n_93480_54040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10113 n_63840_40040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10114 n_91580_40040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10115 n_87020_40040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10116 n_52440_40040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10117 n_90440_40040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10118 n_93480_45640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10119 n_40280_48440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10120 n_79040_40040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10121 n_77140_40040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10122 n_55100_40040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10123 n_40660_45640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10124 n_40660_51240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10125 n_40660_65240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10126 n_41800_68040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10127 n_44840_51240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10128 n_45220_48440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10129 n_54720_42840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10130 n_74860_40040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10131 n_76760_42840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10132 n_41420_48440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10133 n_88920_45640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10134 n_83600_42840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10135 n_51680_42840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10136 n_87020_45640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10137 n_92720_40040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10138 n_63460_42840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10139 n_92340_51240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10140 n_78280_48440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10141 n_64980_48440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10142 n_64600_51240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10143 n_54720_51240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10144 n_63080_51240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10145 n_90440_76440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10146 n_90820_59640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10147 n_91580_79240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10148 n_87400_73640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10149 n_88540_68040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10150 n_89300_54040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10151 n_87780_54040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10152 n_83220_54040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10153 n_91200_54040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10154 n_92340_56840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10155 n_90820_65240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10156 n_88920_70840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10157 n_87400_76440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10158 n_92340_76440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10159 n_83600_84840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10160 n_82080_84840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10161 n_83600_51240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10162 n_80560_51240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10163 n_84740_54040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10164 n_92720_59640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10165 n_90060_79240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10166 n_82080_54040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10167 n_78660_56840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10168 n_83600_56840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10169 n_76380_54040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10170 n_80940_62440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10171 n_76760_56840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10172 n_80560_65240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10173 n_77900_68040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10174 n_76000_70840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10175 n_74860_70840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10176 n_73720_70840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10177 n_75240_76440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10178 n_88920_79240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10179 n_85500_56840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10180 n_87400_48440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10181 n_82080_59640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10182 n_83600_59640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10183 n_82080_65240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10184 n_80560_73640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10185 n_76760_79240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10186 n_80560_79240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10187 n_74860_84840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10188 n_67260_51240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10189 n_70300_51240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10190 n_68780_51240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10191 n_66120_51240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10192 n_79040_51240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10193 n_90820_51240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10194 n_65360_42840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10195 n_92720_42840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10196 n_90440_45640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10197 n_50540_42840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10198 n_85500_42840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10199 n_88920_42840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10200 n_42940_48440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10201 n_76760_45640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10202 n_73340_40040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10203 n_53200_42840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10204 n_44080_48440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10205 n_43320_51240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10206 n_52060_54040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10207 n_59660_62440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10208 n_44840_73640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10209 n_49400_65240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10210 n_61560_62440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10211 n_75240_59640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10212 n_73340_59640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10213 n_55100_56840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10214 n_69160_62440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10215 n_55100_73640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10216 n_50920_70840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10217 n_50920_73640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10218 n_46740_73640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10219 n_40660_76440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10220 n_40660_70840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10221 n_61560_73640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10222 n_58520_73640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10223 n_70300_73640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10224 n_58140_79240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10225 n_54720_68040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10226 n_49400_70840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10227 n_46740_70840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10228 n_63080_73640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10229 n_76760_73640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10230 n_56620_79240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10231 n_61560_79240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10232 n_52060_82040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10233 n_65740_76440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10234 n_44840_76440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10235 n_43320_70840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10236 n_41800_70840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10237 n_40280_82040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10238 n_40280_87640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10239 n_49400_82040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10240 n_54720_84840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10241 n_47120_82040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10242 n_50160_84840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10243 n_70300_76440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10244 n_45220_82040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10245 n_42940_84840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10246 n_40280_84840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10247 n_41420_87640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10248 n_43320_87640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10249 n_46740_84840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10250 n_63080_84840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10251 n_52440_87640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10252 n_59660_84840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10253 n_42940_54040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10254 n_43320_68040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10255 n_43320_76440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10256 n_44080_82040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10257 n_65360_62440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10258 n_66880_62440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10259 n_45220_87640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10260 n_59280_87640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10261 n_51680_84840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10262 n_54340_76440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10263 n_54340_87640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10264 n_64600_84840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10265 n_73340_87640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10266 n_65360_65240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10267 n_67260_65240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10268 n_60040_54040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10269 n_66880_59640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10270 n_70300_65240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10271 n_71820_65240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10272 n_71820_68040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10273 n_70300_68040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10274 n_71820_70840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10275 n_87400_62440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10276 n_88920_62440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10277 n_87020_59640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10278 n_88160_59640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10279 n_85880_62440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10280 n_84740_62440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10281 n_83220_62440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10282 n_85880_73640 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10283 n_83600_76440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10284 n_85500_76440 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10285 n_85500_79240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10286 n_87400_82040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10287 n_83600_82040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10288 n_83600_79240 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10289 n_69920_82040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10290 n_71060_82040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10291 n_72200_82040 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10292 n_44460_56840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10293 n_60040_56840 0 PWL(86000ps 0uA 86030ps 0uA 86031ps 30uA 86059ps 30uA 86060ps 0uA)
I10294 n_90820_68040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10295 n_91200_70840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10296 n_93480_79240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10297 n_87020_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10298 n_93100_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10299 n_90440_62440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10300 n_93100_84840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10301 n_83600_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10302 n_84740_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10303 n_56240_48440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10304 n_61940_48440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10305 n_40660_56840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10306 n_63840_45640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10307 n_79040_42840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10308 n_93480_48440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10309 n_41800_42840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10310 n_48640_40040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10311 n_50920_48440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10312 n_63840_40040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10313 n_88160_40040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10314 n_42940_42840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10315 n_56620_40040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10316 n_67260_40040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10317 n_93480_45640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10318 n_80560_40040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10319 n_40280_40040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10320 n_40280_48440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10321 n_60040_45640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10322 n_77140_40040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10323 n_40660_45640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10324 n_40660_51240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10325 n_42180_73640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10326 n_44460_68040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10327 n_45600_68040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10328 n_43320_62440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10329 n_44460_62440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10330 n_47500_68040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10331 n_46740_65240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10332 n_52060_73640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10333 n_44840_51240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10334 n_45220_48440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10335 n_74860_40040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10336 n_56620_45640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10337 n_41420_48440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10338 n_41420_40040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10339 n_80180_42840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10340 n_88920_45640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10341 n_66880_45640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10342 n_57760_40040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10343 n_44840_45640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10344 n_83600_40040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10345 n_63460_42840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10346 n_51680_48440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10347 n_47880_42840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10348 n_48260_45640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10349 n_90440_48440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10350 n_78280_48440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10351 n_64980_48440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10352 n_41420_54040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10353 n_60040_48440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10354 n_55100_54040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10355 n_81700_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10356 n_80180_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10357 n_90820_84840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10358 n_90820_59640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10359 n_90060_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10360 n_85120_84840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10361 n_91580_79240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10362 n_87400_73640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10363 n_88540_68040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10364 n_87400_65240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10365 n_87400_76440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10366 n_92340_76440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10367 n_82080_84840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10368 n_85880_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10369 n_92720_59640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10370 n_90820_82040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10371 n_77900_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10372 n_79040_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10373 n_78660_56840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10374 n_83600_56840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10375 n_76380_54040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10376 n_80940_62440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10377 n_76760_56840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10378 n_76380_68040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10379 n_78660_65240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10380 n_80560_65240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10381 n_75240_73640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10382 n_73720_79240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10383 n_70300_79240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10384 n_67260_84840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10385 n_65740_84840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10386 n_62320_82040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10387 n_65360_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10388 n_68780_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10389 n_68780_84840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10390 n_70300_84840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10391 n_73720_82040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10392 n_72200_84840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10393 n_86260_54040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10394 n_84740_65240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10395 n_85880_65240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10396 n_87400_68040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10397 n_82080_70840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10398 n_80560_68040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10399 n_77140_70840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10400 n_81700_73640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10401 n_80560_73640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10402 n_78660_73640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10403 n_79040_70840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10404 n_78660_76440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10405 n_78660_79240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10406 n_76760_76440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10407 n_78280_82040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10408 n_76760_84840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10409 n_78660_84840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10410 n_74860_84840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10411 n_76760_82040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10412 n_71820_51240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10413 n_71820_54040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10414 n_68020_54040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10415 n_56620_51240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10416 n_68780_51240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10417 n_59280_51240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10418 n_47880_51240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10419 n_50920_51240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10420 n_41800_56840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10421 n_70300_54040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10422 n_61560_54040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10423 n_66120_51240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10424 n_79040_51240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10425 n_87400_51240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10426 n_49400_48440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10427 n_51680_45640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10428 n_53200_48440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10429 n_65360_42840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10430 n_85500_40040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10431 n_46740_45640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10432 n_61560_40040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10433 n_68020_48440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10434 n_88920_42840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10435 n_82080_42840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10436 n_43320_40040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10437 n_42940_48440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10438 n_53200_45640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10439 n_73340_40040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10440 n_44080_48440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10441 n_43320_51240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10442 n_44840_73640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10443 n_72200_56840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10444 n_49400_65240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10445 n_61560_65240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10446 n_58520_65240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10447 n_59660_68040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10448 n_60420_65240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10449 n_73720_62440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10450 n_66880_68040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10451 n_63080_65240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10452 n_76380_62440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10453 n_75240_59640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10454 n_77520_62440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10455 n_73340_59640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10456 n_61940_68040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10457 n_55100_56840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10458 n_55100_70840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10459 n_53580_70840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10460 n_55100_73640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10461 n_49400_73640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10462 n_55860_68040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10463 n_46740_73640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10464 n_46360_76440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10465 n_40660_76440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10466 n_48260_73640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10467 n_40660_70840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10468 n_49780_76440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10469 n_50920_79240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10470 n_58520_68040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10471 n_58520_73640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10472 n_70300_73640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10473 n_74100_68040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10474 n_75240_68040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10475 n_53580_65240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10476 n_53580_68040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10477 n_54720_68040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10478 n_48260_76440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10479 n_47500_79240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10480 n_48640_79240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10481 n_58520_70840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10482 n_60040_76440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10483 n_60420_70840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10484 n_76760_73640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10485 n_60040_79240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10486 n_63080_79240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10487 n_46360_68040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10488 n_44840_70840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10489 n_44840_76440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10490 n_40660_79240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10491 n_40280_82040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10492 n_43700_79240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10493 n_40280_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10494 n_67260_79240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10495 n_80560_76440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10496 n_50920_82040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10497 n_53580_82040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10498 n_47500_56840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10499 n_44080_59640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10500 n_42940_82040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10501 n_45220_82040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10502 n_40280_84840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10503 n_41420_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10504 n_46740_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10505 n_46740_84840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10506 n_49400_84840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10507 n_52440_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10508 n_49400_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10509 n_64220_82040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10510 n_58140_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10511 n_61940_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10512 n_65360_56840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10513 n_54340_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10514 n_65740_82040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10515 n_53580_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10516 n_56240_76440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10517 n_63460_87640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10518 n_60040_54040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10519 n_70300_59640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10520 n_70300_62440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10521 n_70300_56840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10522 n_70300_70840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10523 n_70300_68040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10524 n_67260_76440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10525 n_65740_79240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10526 n_64600_79240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10527 n_57380_82040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10528 n_55100_79240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10529 n_83220_65240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10530 n_84740_62440 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10531 n_83220_68040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10532 n_83600_70840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10533 n_85500_70840 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10534 n_85880_68040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10535 n_85880_73640 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10536 n_81700_79240 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10537 n_85500_82040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10538 n_68780_82040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10539 n_71060_82040 0 PWL(88000ps 0uA 88030ps 0uA 88031ps 30uA 88059ps 30uA 88060ps 0uA)
I10540 n_93480_79240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10541 n_93100_87640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10542 n_93480_68040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10543 n_93480_76440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10544 n_93100_84840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10545 n_84740_87640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10546 n_65740_40040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10547 n_54720_48440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10548 n_44080_54040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10549 n_40660_56840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10550 n_92340_48440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10551 n_41800_42840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10552 n_50920_48440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10553 n_63840_40040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10554 n_88160_40040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10555 n_67260_40040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10556 n_90440_40040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10557 n_93480_45640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10558 n_80560_40040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10559 n_40280_48440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10560 n_60040_45640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10561 n_82080_48440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10562 n_77140_40040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10563 n_55100_40040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10564 n_40660_45640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10565 n_50160_59640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10566 n_42180_73640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10567 n_44460_68040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10568 n_45600_68040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10569 n_40660_65240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10570 n_41800_68040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10571 n_47500_68040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10572 n_46740_65240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10573 n_52060_73640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10574 n_51300_59640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10575 n_45220_48440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10576 n_54720_42840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10577 n_74860_40040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10578 n_80180_45640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10579 n_56620_45640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10580 n_41420_48440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10581 n_80180_42840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10582 n_88920_45640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10583 n_83600_42840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10584 n_66880_45640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10585 n_83600_40040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10586 n_63460_42840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10587 n_51680_48440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10588 n_48260_45640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10589 n_85120_48440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10590 n_41420_54040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10591 n_49020_51240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10592 n_54720_51240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10593 n_63080_51240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10594 n_81700_87640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10595 n_90820_84840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10596 n_90440_76440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10597 n_92340_65240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10598 n_90060_87640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10599 n_91580_79240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10600 n_92340_76440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10601 n_85880_87640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10602 n_91960_68040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10603 n_90060_79240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10604 n_90820_82040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10605 n_79040_87640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10606 n_76760_65240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10607 n_76380_68040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10608 n_78280_70840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10609 n_75240_73640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10610 n_73720_79240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10611 n_70300_79240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10612 n_67260_84840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10613 n_88920_79240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10614 n_65740_84840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10615 n_62320_82040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10616 n_68780_87640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10617 n_68780_84840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10618 n_71820_87640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10619 n_70300_87640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10620 n_78660_76440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10621 n_78660_79240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10622 n_72200_76440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10623 n_78280_82040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10624 n_76760_84840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10625 n_78660_84840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10626 n_74860_84840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10627 n_67260_51240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10628 n_71820_51240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10629 n_71820_54040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10630 n_70300_51240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10631 n_56620_51240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10632 n_68780_51240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10633 n_59280_51240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10634 n_61940_51240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10635 n_47880_51240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10636 n_41800_56840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10637 n_70300_54040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10638 n_61560_54040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10639 n_83600_48440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10640 n_49400_48440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10641 n_53200_48440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10642 n_65360_42840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10643 n_85500_40040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10644 n_68020_48440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10645 n_85500_42840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10646 n_88920_42840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10647 n_82080_42840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10648 n_42940_48440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10649 n_53200_45640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10650 n_82080_45640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10651 n_73340_40040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10652 n_53200_42840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10653 n_44080_48440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10654 n_57000_54040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10655 n_52060_54040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10656 n_48260_65240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10657 n_59660_62440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10658 n_50920_68040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10659 n_72200_56840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10660 n_53580_59640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10661 n_53580_62440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10662 n_52060_65240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10663 n_49400_65240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10664 n_56620_65240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10665 n_61560_62440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10666 n_61560_65240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10667 n_59660_68040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10668 n_66880_68040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10669 n_63080_65240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10670 n_61940_68040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10671 n_55100_56840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10672 n_69160_62440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10673 n_55100_70840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10674 n_53580_70840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10675 n_50920_70840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10676 n_50920_73640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10677 n_49400_73640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10678 n_55860_68040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10679 n_46360_76440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10680 n_48260_73640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10681 n_49780_76440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10682 n_50920_79240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10683 n_58520_68040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10684 n_61560_73640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10685 n_58140_79240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10686 n_63460_70840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10687 n_65360_70840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10688 n_68780_68040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10689 n_72960_68040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10690 n_55480_48440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10691 n_68780_70840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10692 n_53580_65240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10693 n_53580_68040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10694 n_49400_70840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10695 n_46740_70840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10696 n_48260_76440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10697 n_47500_79240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10698 n_58520_70840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10699 n_60420_70840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10700 n_63080_73640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10701 n_56620_79240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10702 n_60040_79240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10703 n_63080_79240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10704 n_65740_76440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10705 n_58140_51240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10706 n_70300_48440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10707 n_46360_68040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10708 n_44840_70840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10709 n_43320_70840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10710 n_41800_70840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10711 n_40660_79240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10712 n_40280_82040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10713 n_40280_87640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10714 n_57380_76440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10715 n_67260_79240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10716 n_80560_76440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10717 n_50920_82040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10718 n_53580_82040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10719 n_70300_76440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10720 n_40280_84840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10721 n_41420_87640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10722 n_46740_87640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10723 n_46740_84840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10724 n_49400_84840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10725 n_61940_87640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10726 n_42940_54040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10727 n_46740_51240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10728 n_43320_68040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10729 n_43320_76440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10730 n_44080_82040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10731 n_65360_62440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10732 n_66880_62440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10733 n_65360_56840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10734 n_54340_76440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10735 n_56240_76440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10736 n_65360_65240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10737 n_67260_65240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10738 n_66880_59640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10739 n_70300_59640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10740 n_70300_62440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10741 n_70300_56840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10742 n_70300_65240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10743 n_68400_65240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10744 n_71820_68040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10745 n_73720_65240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10746 n_70300_70840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10747 n_67260_76440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10748 n_65740_79240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10749 n_64600_79240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10750 n_57380_82040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10751 n_55100_79240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10752 n_58520_82040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10753 n_59660_82040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10754 n_56240_82040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10755 n_87400_62440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10756 n_87020_59640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10757 n_88160_59640 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10758 n_85880_62440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10759 n_83220_65240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10760 n_83220_68040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10761 n_83600_70840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10762 n_85500_70840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10763 n_85880_68040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10764 n_83600_76440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10765 n_81700_79240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10766 n_85500_76440 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10767 n_85500_79240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10768 n_83600_79240 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10769 n_85500_82040 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10770 n_44460_56840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10771 n_60040_56840 0 PWL(90000ps 0uA 90030ps 0uA 90031ps 30uA 90059ps 30uA 90060ps 0uA)
I10772 n_91200_70840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10773 n_93480_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10774 n_93480_73640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10775 n_93480_76440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10776 n_93100_84840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10777 n_54720_48440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10778 n_56240_48440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10779 n_40280_54040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10780 n_79040_42840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10781 n_93480_48440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10782 n_41800_42840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10783 n_91580_40040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10784 n_87020_40040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10785 n_40660_42840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10786 n_42940_42840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10787 n_67260_40040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10788 n_90440_40040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10789 n_46360_40040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10790 n_40280_40040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10791 n_60040_45640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10792 n_72200_40040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10793 n_79040_40040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10794 n_82080_48440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10795 n_77140_40040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10796 n_50160_59640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10797 n_42180_73640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10798 n_44460_68040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10799 n_45600_68040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10800 n_40660_65240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10801 n_41800_68040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10802 n_47500_68040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10803 n_46740_65240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10804 n_52060_73640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10805 n_51300_59640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10806 n_74860_40040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10807 n_80180_45640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10808 n_76760_42840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10809 n_71820_42840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10810 n_56620_45640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10811 n_41420_40040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10812 n_49400_40040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10813 n_83600_42840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10814 n_66880_45640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10815 n_44840_45640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10816 n_43700_42840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10817 n_87020_45640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10818 n_92720_40040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10819 n_48260_45640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10820 n_90440_48440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10821 n_78280_48440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10822 n_47880_54040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10823 n_55100_54040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10824 n_54720_51240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10825 n_90820_84840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10826 n_90440_76440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10827 n_90440_73640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10828 n_91580_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10829 n_87400_73640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10830 n_87400_76440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10831 n_92340_76440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10832 n_92340_73640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10833 n_90060_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10834 n_90820_82040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10835 n_80940_62440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10836 n_76760_56840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10837 n_79040_68040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10838 n_75240_73640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10839 n_74860_70840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10840 n_73720_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10841 n_70300_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10842 n_67260_84840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10843 n_71820_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10844 n_88920_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10845 n_65740_84840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10846 n_62320_82040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10847 n_68780_84840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10848 n_84740_65240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10849 n_82080_68040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10850 n_80560_68040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10851 n_77140_70840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10852 n_80560_73640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10853 n_81700_76440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10854 n_79040_70840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10855 n_78660_76440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10856 n_78660_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10857 n_78280_82040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10858 n_76760_84840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10859 n_78660_84840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10860 n_70300_51240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10861 n_68020_54040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10862 n_49780_54040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10863 n_79040_51240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10864 n_87400_51240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10865 n_49400_48440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10866 n_92720_42840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10867 n_90440_45640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10868 n_45220_42840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10869 n_46740_45640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10870 n_68020_48440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10871 n_85500_42840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10872 n_51300_40040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10873 n_43320_40040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10874 n_53200_45640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10875 n_73720_45640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10876 n_76760_45640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10877 n_82080_45640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10878 n_73340_40040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10879 n_58900_48440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10880 n_57000_54040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10881 n_48260_65240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10882 n_59660_62440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10883 n_50920_68040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10884 n_72200_56840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10885 n_53580_59640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10886 n_53580_62440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10887 n_52060_65240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10888 n_49400_65240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10889 n_56620_65240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10890 n_61560_62440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10891 n_61560_65240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10892 n_59660_68040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10893 n_60800_68040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10894 n_60040_73640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10895 n_63080_65240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10896 n_76380_59640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10897 n_61940_68040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10898 n_59660_70840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10899 n_55100_56840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10900 n_69160_62440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10901 n_55100_70840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10902 n_53580_70840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10903 n_50920_70840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10904 n_50920_73640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10905 n_49400_73640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10906 n_55860_68040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10907 n_46360_76440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10908 n_48260_73640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10909 n_49780_76440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10910 n_50920_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10911 n_58520_73640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10912 n_70300_73640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10913 n_66880_73640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10914 n_58140_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10915 n_55480_48440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10916 n_53580_65240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10917 n_53580_68040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10918 n_49400_70840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10919 n_46740_70840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10920 n_48260_76440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10921 n_47500_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10922 n_58520_70840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10923 n_60420_70840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10924 n_76760_73640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10925 n_56620_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10926 n_60040_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10927 n_63080_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10928 n_65740_76440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10929 n_68400_73640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10930 n_58140_51240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10931 n_70300_48440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10932 n_46360_68040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10933 n_44840_70840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10934 n_43320_70840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10935 n_41800_70840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10936 n_40660_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10937 n_40280_82040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10938 n_40280_87640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10939 n_57380_76440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10940 n_67260_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10941 n_80560_76440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10942 n_50920_82040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10943 n_53580_82040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10944 n_70300_76440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10945 n_52820_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10946 n_40280_84840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10947 n_41420_87640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10948 n_46740_87640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10949 n_46740_84840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10950 n_49400_84840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10951 n_61940_87640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10952 n_46740_51240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10953 n_43320_68040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10954 n_43320_76440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10955 n_44080_82040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10956 n_65360_62440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10957 n_66880_62440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10958 n_65360_56840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10959 n_68780_56840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10960 n_54340_76440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10961 n_65360_65240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10962 n_67260_65240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10963 n_67260_56840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10964 n_66880_59640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10965 n_70300_59640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10966 n_70300_56840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10967 n_70300_65240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10968 n_68400_65240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10969 n_71820_68040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10970 n_70300_70840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10971 n_70300_68040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10972 n_67260_76440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10973 n_65740_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10974 n_64600_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10975 n_53960_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10976 n_64600_76440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10977 n_55100_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10978 n_56240_82040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10979 n_87400_62440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10980 n_87020_59640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10981 n_88160_59640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10982 n_85880_62440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10983 n_83220_65240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10984 n_83220_68040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10985 n_83600_70840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10986 n_83220_73640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10987 n_85880_73640 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10988 n_83600_76440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10989 n_81700_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10990 n_85500_76440 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10991 n_85500_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10992 n_83600_79240 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10993 n_85500_82040 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10994 n_44460_56840 0 PWL(92000ps 0uA 92030ps 0uA 92031ps 30uA 92059ps 30uA 92060ps 0uA)
I10995 n_91200_70840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I10996 n_91960_87640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I10997 n_93480_76440 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I10998 n_93100_84840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I10999 n_84740_87640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11000 n_54720_48440 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11001 n_61940_48440 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11002 n_44080_54040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11003 n_93480_48440 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11004 n_48640_40040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11005 n_70300_40040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11006 n_91580_40040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11007 n_87020_40040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11008 n_52440_40040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11009 n_40660_42840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11010 n_42940_42840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11011 n_67260_40040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11012 n_80560_40040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11013 n_40280_48440 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11014 n_60040_45640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11015 n_72200_40040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11016 n_79040_40040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11017 n_55100_40040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11018 n_40660_45640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11019 n_40660_51240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11020 n_44840_51240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11021 n_45220_48440 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11022 n_54720_42840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11023 n_76760_42840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11024 n_71820_42840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11025 n_56620_45640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11026 n_41420_48440 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11027 n_80180_42840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11028 n_66880_45640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11029 n_44840_45640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11030 n_43700_42840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11031 n_51680_42840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11032 n_87020_45640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11033 n_92720_40040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11034 n_68400_40040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11035 n_47880_42840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11036 n_90440_48440 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11037 n_49020_51240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11038 n_60040_48440 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11039 n_54720_51240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11040 n_81700_87640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11041 n_90820_84840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11042 n_90440_76440 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11043 n_87400_84840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11044 n_87400_73640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11045 n_87400_76440 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11046 n_88920_82040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11047 n_87400_56840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11048 n_90820_56840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11049 n_77520_54040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11050 n_87400_79240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11051 n_89300_73640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11052 n_92340_73640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11053 n_88920_76440 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11054 n_89300_84840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11055 n_80560_84840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11056 n_77900_87640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11057 n_79040_87640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11058 n_79040_54040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11059 n_80560_54040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11060 n_80560_56840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11061 n_82080_56840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11062 n_78660_56840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11063 n_76760_65240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11064 n_78660_65240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11065 n_77900_68040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11066 n_76000_70840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11067 n_79040_68040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11068 n_75240_73640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11069 n_73720_79240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11070 n_70300_79240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11071 n_67260_84840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11072 n_71820_79240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11073 n_88920_79240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11074 n_65740_84840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11075 n_65360_87640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11076 n_73720_82040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11077 n_85500_59640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11078 n_84740_65240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11079 n_82080_68040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11080 n_80560_68040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11081 n_77140_70840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11082 n_80560_73640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11083 n_79040_70840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11084 n_80560_79240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11085 n_80180_82040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11086 n_76760_84840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11087 n_78660_84840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11088 n_60800_51240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11089 n_67260_51240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11090 n_71820_51240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11091 n_71820_54040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11092 n_53200_51240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11093 n_53580_54040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11094 n_68020_54040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11095 n_56620_51240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11096 n_68780_51240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11097 n_61940_51240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11098 n_46360_54040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11099 n_49780_54040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11100 n_47880_51240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11101 n_70300_54040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11102 n_61560_54040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11103 n_87400_51240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11104 n_51680_45640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11105 n_70300_42840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11106 n_92720_42840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11107 n_90440_45640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11108 n_50540_42840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11109 n_45220_42840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11110 n_46740_45640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11111 n_68020_48440 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11112 n_82080_42840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11113 n_42940_48440 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11114 n_53200_45640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11115 n_73720_45640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11116 n_76760_45640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11117 n_53200_42840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11118 n_44080_48440 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11119 n_43320_51240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11120 n_57000_54040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11121 n_72200_56840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11122 n_55100_56840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11123 n_70300_73640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11124 n_56620_73640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11125 n_58140_79240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11126 n_68780_70840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11127 n_63080_73640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11128 n_76760_73640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11129 n_56620_79240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11130 n_60040_79240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11131 n_61560_79240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11132 n_52060_82040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11133 n_65740_76440 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11134 n_58140_51240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11135 n_50920_82040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11136 n_49400_82040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11137 n_54720_84840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11138 n_53580_82040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11139 n_70300_76440 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11140 n_47500_56840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11141 n_46740_84840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11142 n_63080_84840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11143 n_49400_84840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11144 n_61940_87640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11145 n_42940_54040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11146 n_46740_51240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11147 n_68780_56840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11148 n_67260_56840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11149 n_66880_59640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11150 n_70300_59640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11151 n_70300_56840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11152 n_73720_65240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11153 n_70300_68040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11154 n_59660_82040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11155 n_56240_82040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11156 n_85500_70840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11157 n_83220_73640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11158 n_84740_73640 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11159 n_83600_76440 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11160 n_81700_79240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11161 n_85500_76440 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11162 n_87400_82040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11163 n_85500_82040 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11164 n_43320_65240 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11165 n_60040_56840 0 PWL(94000ps 0uA 94030ps 0uA 94031ps 30uA 94059ps 30uA 94060ps 0uA)
I11166 n_93480_79240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11167 n_93100_87640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11168 n_93480_76440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11169 n_54720_48440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11170 n_65740_45640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11171 n_40280_54040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11172 n_44080_54040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11173 n_40660_56840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11174 n_93480_48440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11175 n_93480_54040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11176 n_92340_48440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11177 n_41800_42840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11178 n_48640_40040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11179 n_50920_48440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11180 n_91580_40040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11181 n_87020_40040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11182 n_88160_40040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11183 n_52440_40040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11184 n_40660_42840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11185 n_42940_42840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11186 n_56620_40040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11187 n_80560_40040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11188 n_40280_40040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11189 n_60040_45640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11190 n_82080_48440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11191 n_40660_45640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11192 n_40660_51240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11193 n_44840_51240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11194 n_45220_48440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11195 n_80180_45640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11196 n_56620_45640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11197 n_41420_40040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11198 n_80180_42840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11199 n_57760_40040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11200 n_44840_45640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11201 n_43700_42840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11202 n_51680_42840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11203 n_83600_40040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11204 n_87020_45640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11205 n_92720_40040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11206 n_51680_48440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11207 n_47880_42840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11208 n_48260_45640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11209 n_85120_48440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11210 n_92340_51240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11211 n_90440_48440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11212 n_41420_54040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11213 n_49020_51240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11214 n_47880_54040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11215 n_64600_51240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11216 n_54720_51240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11217 n_90440_76440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11218 n_90060_87640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11219 n_91580_79240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11220 n_92340_76440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11221 n_85880_87640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11222 n_87400_56840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11223 n_90820_56840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11224 n_77520_54040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11225 n_87400_79240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11226 n_89300_73640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11227 n_92340_73640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11228 n_88920_76440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11229 n_89300_84840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11230 n_90820_82040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11231 n_80560_84840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11232 n_77900_87640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11233 n_79040_54040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11234 n_80560_54040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11235 n_80560_56840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11236 n_82080_56840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11237 n_78660_56840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11238 n_76760_65240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11239 n_78660_65240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11240 n_77900_68040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11241 n_79040_68040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11242 n_73720_70840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11243 n_73720_73640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11244 n_88920_79240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11245 n_62320_82040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11246 n_65360_87640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11247 n_68780_84840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11248 n_71820_87640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11249 n_70300_87640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11250 n_73720_82040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11251 n_82080_70840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11252 n_80560_68040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11253 n_77140_70840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11254 n_81700_73640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11255 n_81700_76440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11256 n_78660_73640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11257 n_79040_70840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11258 n_78660_76440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11259 n_78660_79240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11260 n_76760_76440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11261 n_72200_76440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11262 n_78280_82040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11263 n_76760_79240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11264 n_80180_82040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11265 n_74860_84840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11266 n_60800_51240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11267 n_67260_51240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11268 n_71820_51240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11269 n_71820_54040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11270 n_53200_51240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11271 n_53580_54040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11272 n_68020_54040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11273 n_56620_51240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11274 n_46360_54040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11275 n_47880_51240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11276 n_52060_51240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11277 n_70300_54040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11278 n_61560_54040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11279 n_87400_51240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11280 n_90820_51240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11281 n_83600_48440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11282 n_49400_48440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11283 n_51680_45640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11284 n_53200_48440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11285 n_92720_42840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11286 n_90440_45640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11287 n_85500_40040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11288 n_50540_42840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11289 n_45220_42840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11290 n_46740_45640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11291 n_61560_40040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11292 n_82080_42840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11293 n_43320_40040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11294 n_53200_45640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11295 n_82080_45640 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11296 n_44080_48440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11297 n_43320_51240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11298 n_52060_54040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11299 n_55480_48440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11300 n_63080_79240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11301 n_61560_79240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11302 n_65740_76440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11303 n_70300_48440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11304 n_57380_76440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11305 n_67260_79240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11306 n_80560_76440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11307 n_70300_76440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11308 n_46740_51240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11309 n_65360_56840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11310 n_70300_70840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11311 n_70300_68040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11312 n_71820_70840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11313 n_67260_76440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11314 n_68780_76440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11315 n_65740_79240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11316 n_64600_79240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11317 n_53960_79240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11318 n_64600_76440 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11319 n_59660_82040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11320 n_56240_82040 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11321 n_43320_65240 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11322 n_44460_56840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11323 n_60040_56840 0 PWL(96000ps 0uA 96030ps 0uA 96031ps 30uA 96059ps 30uA 96060ps 0uA)
I11324 n_93480_79240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11325 n_87020_87640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11326 n_93100_87640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11327 n_93480_73640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11328 n_93100_84840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11329 n_84740_87640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11330 n_56240_48440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11331 n_44080_54040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11332 n_93480_48440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11333 n_48640_40040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11334 n_63840_40040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11335 n_70300_40040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11336 n_91580_40040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11337 n_40660_42840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11338 n_42940_42840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11339 n_56620_40040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11340 n_60040_45640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11341 n_72200_40040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11342 n_79040_40040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11343 n_55100_40040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11344 n_40660_45640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11345 n_40660_51240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11346 n_43320_59640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11347 n_40660_65240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11348 n_41800_68040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11349 n_46740_59640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11350 n_44840_51240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11351 n_45220_48440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11352 n_54720_42840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11353 n_76760_42840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11354 n_71820_42840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11355 n_56620_45640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11356 n_57760_40040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11357 n_44840_45640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11358 n_43700_42840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11359 n_92720_40040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11360 n_68400_40040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11361 n_63460_42840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11362 n_47880_42840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11363 n_90440_48440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11364 n_49020_51240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11365 n_55100_54040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11366 n_81700_87640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11367 n_90820_84840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11368 n_90440_73640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11369 n_90060_87640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11370 n_85120_84840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11371 n_91580_79240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11372 n_92340_76440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11373 n_82080_84840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11374 n_85880_87640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11375 n_87400_56840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11376 n_90820_56840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11377 n_77520_54040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11378 n_87400_79240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11379 n_92340_73640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11380 n_90820_82040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11381 n_80560_84840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11382 n_77900_87640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11383 n_81700_82040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11384 n_79040_54040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11385 n_80560_54040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11386 n_80560_56840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11387 n_82080_56840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11388 n_78660_56840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11389 n_76760_65240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11390 n_78660_65240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11391 n_77900_68040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11392 n_79040_68040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11393 n_75240_76440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11394 n_70300_79240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11395 n_67260_84840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11396 n_88920_79240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11397 n_67260_87640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11398 n_65360_87640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11399 n_68780_87640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11400 n_68780_84840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11401 n_70300_84840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11402 n_73720_82040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11403 n_72200_84840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11404 n_80560_68040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11405 n_77140_70840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11406 n_76760_76440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11407 n_78280_82040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11408 n_76760_84840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11409 n_76380_87640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11410 n_74860_84840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11411 n_76760_82040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11412 n_68020_54040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11413 n_50920_51240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11414 n_87400_51240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11415 n_51680_45640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11416 n_65360_42840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11417 n_70300_42840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11418 n_92720_42840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11419 n_45220_42840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11420 n_46740_45640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11421 n_61560_40040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11422 n_53200_45640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11423 n_73720_45640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11424 n_76760_45640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11425 n_53200_42840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11426 n_44080_48440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11427 n_43320_51240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11428 n_58900_48440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11429 n_49780_56840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11430 n_48260_62440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11431 n_52060_54040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11432 n_48260_65240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11433 n_49780_62440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11434 n_59660_62440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11435 n_44840_73640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11436 n_50920_68040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11437 n_72200_56840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11438 n_56620_65240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11439 n_61560_62440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11440 n_61560_65240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11441 n_59660_68040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11442 n_60800_68040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11443 n_60040_73640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11444 n_63080_65240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11445 n_61940_68040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11446 n_59660_70840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11447 n_49400_73640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11448 n_55860_68040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11449 n_46740_73640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11450 n_46360_76440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11451 n_40660_76440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11452 n_48260_73640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11453 n_40660_70840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11454 n_49780_76440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11455 n_50920_79240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11456 n_58520_73640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11457 n_56620_73640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11458 n_58140_79240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11459 n_68780_70840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11460 n_48260_76440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11461 n_47500_79240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11462 n_48640_79240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11463 n_58520_70840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11464 n_60040_76440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11465 n_60420_70840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11466 n_63080_73640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11467 n_60040_79240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11468 n_63080_79240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11469 n_52060_82040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11470 n_65740_76440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11471 n_40660_79240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11472 n_40280_82040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11473 n_43700_79240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11474 n_40280_87640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11475 n_67260_79240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11476 n_80560_76440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11477 n_50920_82040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11478 n_53580_82040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11479 n_70300_76440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11480 n_52820_79240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11481 n_40280_84840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11482 n_41420_87640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11483 n_46740_87640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11484 n_46740_84840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11485 n_49400_84840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11486 n_52440_87640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11487 n_49400_87640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11488 n_64220_82040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11489 n_58140_87640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11490 n_61940_87640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11491 n_46740_51240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11492 n_43320_68040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11493 n_43320_76440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11494 n_44080_82040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11495 n_65360_62440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11496 n_66880_62440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11497 n_54340_87640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11498 n_65740_82040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11499 n_53580_87640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11500 n_56240_76440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11501 n_63460_87640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11502 n_65360_65240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11503 n_67260_65240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11504 n_60040_54040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11505 n_71820_59640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11506 n_70300_65240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11507 n_71820_65240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11508 n_71820_68040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11509 n_70300_68040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11510 n_71820_70840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11511 n_55100_79240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11512 n_58520_82040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11513 n_59660_82040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11514 n_56620_84840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11515 n_87400_62440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11516 n_87020_59640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11517 n_88160_59640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11518 n_85880_62440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11519 n_83220_65240 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11520 n_83220_68040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11521 n_83600_70840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11522 n_85500_70840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11523 n_84740_73640 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11524 n_83600_76440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11525 n_85500_76440 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11526 n_87400_82040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11527 n_68780_82040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11528 n_71060_82040 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11529 n_44460_56840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11530 n_60040_56840 0 PWL(98000ps 0uA 98030ps 0uA 98031ps 30uA 98059ps 30uA 98060ps 0uA)
I11531 n_93480_79240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11532 n_91960_87640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11533 n_93100_87640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11534 n_93480_73640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11535 n_93100_84840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11536 n_84740_87640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11537 n_65740_45640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11538 n_40280_54040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11539 n_93480_54040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11540 n_41800_42840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11541 n_63840_40040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11542 n_87020_40040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11543 n_42940_42840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11544 n_80560_40040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11545 n_79040_40040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11546 n_82080_48440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11547 n_43320_59640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11548 n_46740_59640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11549 n_80180_45640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11550 n_76760_42840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11551 n_80180_42840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11552 n_44840_45640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11553 n_87020_45640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11554 n_63460_42840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11555 n_48260_45640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11556 n_92340_51240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11557 n_47880_54040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11558 n_64600_51240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11559 n_81700_87640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11560 n_90820_84840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11561 n_90440_73640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11562 n_90060_87640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11563 n_87400_84840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11564 n_91580_79240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11565 n_92340_76440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11566 n_88920_82040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11567 n_85880_87640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11568 n_87400_56840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11569 n_90820_56840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11570 n_77520_54040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11571 n_87400_79240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11572 n_92340_73640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11573 n_90820_82040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11574 n_80560_84840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11575 n_77900_87640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11576 n_81700_82040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11577 n_79040_54040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11578 n_80560_54040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11579 n_80560_56840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11580 n_82080_56840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11581 n_78660_56840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11582 n_76760_65240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11583 n_78660_65240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11584 n_77900_68040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11585 n_76000_70840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11586 n_75240_73640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11587 n_73720_70840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11588 n_75240_76440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11589 n_73720_79240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11590 n_73720_73640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11591 n_88920_79240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11592 n_62320_82040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11593 n_70300_84840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11594 n_72200_84840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11595 n_82080_70840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11596 n_81700_73640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11597 n_78660_73640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11598 n_79040_70840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11599 n_78660_79240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11600 n_76760_76440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11601 n_76760_79240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11602 n_80560_79240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11603 n_78660_84840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11604 n_76380_87640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11605 n_74860_84840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11606 n_68780_51240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11607 n_49780_54040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11608 n_90820_51240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11609 n_49400_48440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11610 n_65360_42840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11611 n_90440_45640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11612 n_46740_45640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11613 n_82080_42840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11614 n_76760_45640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11615 n_82080_45640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11616 n_49780_56840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11617 n_48260_62440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11618 n_48260_65240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11619 n_49780_62440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11620 n_59660_62440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11621 n_44840_73640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11622 n_50920_68040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11623 n_72200_56840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11624 n_56620_65240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11625 n_61560_62440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11626 n_61560_65240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11627 n_59660_68040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11628 n_60800_68040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11629 n_60040_73640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11630 n_63080_65240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11631 n_61940_68040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11632 n_59660_70840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11633 n_55100_56840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11634 n_69160_62440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11635 n_49400_73640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11636 n_55860_68040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11637 n_46740_73640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11638 n_46360_76440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11639 n_40660_76440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11640 n_48260_73640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11641 n_40660_70840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11642 n_49780_76440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11643 n_50920_79240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11644 n_58520_73640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11645 n_56620_73640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11646 n_58140_79240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11647 n_55480_48440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11648 n_48260_76440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11649 n_47500_79240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11650 n_48640_79240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11651 n_58520_70840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11652 n_60040_76440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11653 n_60420_70840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11654 n_63080_73640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11655 n_60040_79240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11656 n_63080_79240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11657 n_52060_82040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11658 n_65740_76440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11659 n_40660_79240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11660 n_40280_82040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11661 n_43700_79240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11662 n_44080_84840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11663 n_40280_87640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11664 n_67260_79240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11665 n_80560_76440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11666 n_50920_82040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11667 n_54720_84840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11668 n_47120_82040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11669 n_53580_82040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11670 n_50160_84840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11671 n_70300_76440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11672 n_41420_87640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11673 n_46740_87640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11674 n_63080_84840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11675 n_49400_84840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11676 n_52440_87640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11677 n_58140_87640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11678 n_61940_87640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11679 n_42940_54040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11680 n_65360_62440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11681 n_66880_62440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11682 n_45220_87640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11683 n_51680_84840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11684 n_54340_87640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11685 n_53580_87640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11686 n_56240_76440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11687 n_63460_87640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11688 n_65360_65240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11689 n_67260_65240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11690 n_68400_65240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11691 n_71820_65240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11692 n_73720_65240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11693 n_55100_79240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11694 n_58520_82040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11695 n_56240_82040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11696 n_56620_84840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11697 n_87400_62440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11698 n_87020_59640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11699 n_88160_59640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11700 n_85880_62440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11701 n_83220_65240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11702 n_83220_68040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11703 n_83600_70840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11704 n_85500_70840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11705 n_84740_73640 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11706 n_83600_76440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11707 n_85500_76440 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11708 n_85500_79240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11709 n_83600_82040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11710 n_69920_82040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11711 n_71060_82040 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11712 n_43320_65240 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11713 n_44460_56840 0 PWL(100000ps 0uA 100030ps 0uA 100031ps 30uA 100059ps 30uA 100060ps 0uA)
I11714 n_91960_87640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11715 n_93100_84840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11716 n_54720_48440 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11717 n_56240_48440 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11718 n_61940_48440 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11719 n_40280_54040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11720 n_44080_54040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11721 n_79040_42840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11722 n_93480_48440 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11723 n_92340_48440 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11724 n_41800_42840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11725 n_48640_40040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11726 n_91580_40040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11727 n_87020_40040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11728 n_88160_40040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11729 n_52440_40040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11730 n_42940_42840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11731 n_56620_40040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11732 n_67260_40040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11733 n_90440_40040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11734 n_93480_45640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11735 n_80560_40040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11736 n_46360_40040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11737 n_40280_40040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11738 n_60040_45640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11739 n_79040_40040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11740 n_82080_48440 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11741 n_80180_45640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11742 n_76760_42840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11743 n_56620_45640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11744 n_41420_40040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11745 n_49400_40040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11746 n_80180_42840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11747 n_88920_45640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11748 n_83600_42840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11749 n_66880_45640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11750 n_57760_40040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11751 n_44840_45640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11752 n_51680_42840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11753 n_83600_40040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11754 n_87020_45640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11755 n_92720_40040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11756 n_47880_42840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11757 n_48260_45640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11758 n_85120_48440 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11759 n_90440_48440 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11760 n_78280_48440 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11761 n_49020_51240 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11762 n_47880_54040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11763 n_60040_48440 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11764 n_55100_54040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11765 n_54720_51240 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11766 n_90820_84840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11767 n_87400_84840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11768 n_88920_82040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11769 n_90820_82040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11770 n_80940_62440 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11771 n_76760_56840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11772 n_79040_68040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11773 n_67260_84840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11774 n_71820_79240 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11775 n_67260_87640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11776 n_62320_82040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11777 n_65360_87640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11778 n_73720_82040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11779 n_85500_56840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11780 n_82080_59640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11781 n_85500_59640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11782 n_84740_65240 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11783 n_83600_59640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11784 n_82080_68040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11785 n_80560_68040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11786 n_77140_70840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11787 n_78660_79240 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11788 n_76760_76440 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11789 n_72200_76440 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11790 n_78280_82040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11791 n_76760_79240 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11792 n_80560_79240 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11793 n_76760_84840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11794 n_78660_84840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11795 n_74860_82040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11796 n_70300_51240 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11797 n_68020_54040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11798 n_61940_51240 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11799 n_49780_54040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11800 n_50920_51240 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11801 n_79040_51240 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11802 n_87400_51240 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11803 n_83600_48440 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11804 n_49400_48440 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11805 n_51680_45640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11806 n_92720_42840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11807 n_90440_45640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11808 n_85500_40040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11809 n_50540_42840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11810 n_46740_45640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11811 n_61560_40040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11812 n_68020_48440 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11813 n_85500_42840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11814 n_88920_42840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11815 n_82080_42840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11816 n_51300_40040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11817 n_43320_40040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11818 n_53200_45640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11819 n_76760_45640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11820 n_82080_45640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11821 n_72200_56840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11822 n_76380_59640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11823 n_55100_56840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11824 n_69160_62440 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11825 n_68780_70840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11826 n_58140_51240 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11827 n_54720_84840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11828 n_47120_82040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11829 n_53580_82040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11830 n_47500_56840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11831 n_46740_84840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11832 n_63080_84840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11833 n_49400_84840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11834 n_61940_87640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11835 n_42940_54040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11836 n_60040_54040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11837 n_66880_59640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11838 n_70300_59640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11839 n_70300_62440 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11840 n_70300_56840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11841 n_71820_59640 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11842 n_70300_65240 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11843 n_68400_65240 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11844 n_71820_68040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11845 n_73720_65240 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11846 n_70300_68040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11847 n_68780_76440 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11848 n_55100_79240 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11849 n_59660_82040 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11850 n_43320_65240 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11851 n_60040_56840 0 PWL(102000ps 0uA 102030ps 0uA 102031ps 30uA 102059ps 30uA 102060ps 0uA)
I11852 n_91960_87640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11853 n_87020_87640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11854 n_93100_84840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11855 n_54720_48440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11856 n_65740_45640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11857 n_61940_48440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11858 n_40280_54040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11859 n_44080_54040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11860 n_40660_56840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11861 n_79040_42840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11862 n_93480_54040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11863 n_92340_48440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11864 n_41800_42840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11865 n_48640_40040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11866 n_50920_48440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11867 n_88160_40040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11868 n_52440_40040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11869 n_40660_42840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11870 n_67260_40040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11871 n_93480_45640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11872 n_80560_40040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11873 n_40280_40040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11874 n_40280_48440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11875 n_72200_40040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11876 n_55100_40040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11877 n_40660_45640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11878 n_43320_59640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11879 n_46740_59640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11880 n_45220_48440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11881 n_54720_42840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11882 n_71820_42840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11883 n_41420_48440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11884 n_41420_40040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11885 n_80180_42840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11886 n_88920_45640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11887 n_66880_45640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11888 n_43700_42840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11889 n_51680_42840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11890 n_83600_40040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11891 n_51680_48440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11892 n_47880_42840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11893 n_48260_45640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11894 n_85120_48440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11895 n_92340_51240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11896 n_78280_48440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11897 n_41420_54040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11898 n_49020_51240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11899 n_47880_54040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11900 n_60040_48440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11901 n_64600_51240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11902 n_54720_51240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11903 n_90820_84840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11904 n_85120_84840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11905 n_87400_84840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11906 n_88920_82040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11907 n_82080_84840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11908 n_90820_82040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11909 n_80940_62440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11910 n_76760_56840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11911 n_76000_70840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11912 n_75240_73640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11913 n_73720_70840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11914 n_73720_79240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11915 n_73720_73640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11916 n_67260_84840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11917 n_71820_79240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11918 n_67260_87640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11919 n_62320_82040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11920 n_65360_87640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11921 n_70300_87640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11922 n_73720_82040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11923 n_85500_56840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11924 n_82080_59640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11925 n_85500_59640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11926 n_84740_65240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11927 n_83600_59640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11928 n_82080_68040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11929 n_82080_70840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11930 n_81700_73640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11931 n_78660_73640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11932 n_79040_70840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11933 n_78660_79240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11934 n_76760_76440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11935 n_72200_76440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11936 n_78280_82040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11937 n_76760_79240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11938 n_80560_79240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11939 n_80180_82040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11940 n_76760_84840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11941 n_78660_84840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11942 n_74860_82040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11943 n_76760_82040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11944 n_70300_51240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11945 n_68780_51240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11946 n_61940_51240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11947 n_49780_54040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11948 n_50920_51240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11949 n_52060_51240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11950 n_79040_51240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11951 n_90820_51240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11952 n_83600_48440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11953 n_49400_48440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11954 n_51680_45640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11955 n_53200_48440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11956 n_85500_40040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11957 n_50540_42840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11958 n_45220_42840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11959 n_68020_48440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11960 n_88920_42840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11961 n_82080_42840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11962 n_43320_40040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11963 n_42940_48440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11964 n_73720_45640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11965 n_53200_42840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11966 n_44080_48440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11967 n_49780_56840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11968 n_48260_62440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11969 n_52060_54040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11970 n_48260_65240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11971 n_49780_62440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11972 n_59660_62440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11973 n_44840_73640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11974 n_50920_68040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11975 n_72200_56840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11976 n_56620_65240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11977 n_61560_62440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11978 n_61560_65240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11979 n_59660_68040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11980 n_60800_68040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11981 n_60040_73640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11982 n_63080_65240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11983 n_76380_59640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11984 n_61940_68040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11985 n_59660_70840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11986 n_55100_56840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11987 n_49400_73640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11988 n_55860_68040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11989 n_46740_73640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11990 n_46360_76440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11991 n_40660_76440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11992 n_48260_73640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11993 n_40660_70840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11994 n_49780_76440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11995 n_50920_79240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11996 n_58520_73640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11997 n_56620_73640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11998 n_58140_79240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I11999 n_68780_70840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12000 n_48260_76440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12001 n_47500_79240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12002 n_48640_79240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12003 n_58520_70840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12004 n_60040_76440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12005 n_60420_70840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12006 n_63080_73640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12007 n_56620_79240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12008 n_52060_82040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12009 n_58140_51240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12010 n_70300_48440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12011 n_40660_79240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12012 n_40280_82040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12013 n_43700_79240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12014 n_44080_84840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12015 n_40280_87640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12016 n_57380_76440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12017 n_49400_82040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12018 n_54720_84840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12019 n_53580_82040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12020 n_50160_84840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12021 n_47500_56840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12022 n_41420_87640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12023 n_46740_87640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12024 n_63080_84840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12025 n_49400_84840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12026 n_49400_87640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12027 n_64220_82040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12028 n_61940_87640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12029 n_65360_62440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12030 n_66880_62440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12031 n_45220_87640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12032 n_51680_84840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12033 n_65740_82040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12034 n_65360_65240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12035 n_67260_65240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12036 n_66880_59640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12037 n_70300_59640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12038 n_70300_62440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12039 n_70300_56840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12040 n_55100_79240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12041 n_59660_82040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12042 n_87400_62440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12043 n_87020_59640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12044 n_88160_59640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12045 n_85880_62440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12046 n_83220_65240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12047 n_83220_68040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12048 n_83600_70840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12049 n_85500_70840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12050 n_84740_73640 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12051 n_83600_76440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12052 n_85500_76440 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12053 n_85500_79240 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12054 n_83600_82040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12055 n_69920_82040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12056 n_68780_82040 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12057 n_44460_56840 0 PWL(104000ps 0uA 104030ps 0uA 104031ps 30uA 104059ps 30uA 104060ps 0uA)
I12058 n_90820_68040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12059 n_93480_79240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12060 n_93480_56840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12061 n_90440_62440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12062 n_93100_84840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12063 n_83600_87640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12064 n_65740_40040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12065 n_54720_48440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12066 n_56240_48440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12067 n_40280_54040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12068 n_44080_54040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12069 n_40660_56840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12070 n_63840_45640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12071 n_79040_42840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12072 n_93480_48440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12073 n_41800_42840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12074 n_48640_40040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12075 n_50920_48440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12076 n_63840_40040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12077 n_70300_40040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12078 n_91580_40040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12079 n_52440_40040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12080 n_40660_42840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12081 n_42940_42840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12082 n_56620_40040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12083 n_90440_40040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12084 n_40280_48440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12085 n_60040_45640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12086 n_72200_40040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12087 n_77140_40040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12088 n_55100_40040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12089 n_40660_45640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12090 n_43320_59640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12091 n_40660_65240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12092 n_41800_68040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12093 n_46740_59640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12094 n_45220_48440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12095 n_54720_42840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12096 n_74860_40040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12097 n_71820_42840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12098 n_56620_45640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12099 n_41420_48440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12100 n_83600_42840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12101 n_57760_40040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12102 n_44840_45640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12103 n_43700_42840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12104 n_51680_42840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12105 n_92720_40040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12106 n_68400_40040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12107 n_63460_42840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12108 n_51680_48440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12109 n_47880_42840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12110 n_48260_45640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12111 n_90440_48440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12112 n_78280_48440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12113 n_64980_48440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12114 n_41420_54040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12115 n_49020_51240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12116 n_47880_54040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12117 n_55100_54040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12118 n_54720_51240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12119 n_63080_51240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12120 n_80180_87640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12121 n_90820_84840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12122 n_90820_59640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12123 n_88920_56840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12124 n_91580_79240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12125 n_88540_68040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12126 n_68780_79240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12127 n_83220_54040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12128 n_91200_54040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12129 n_92340_56840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12130 n_90820_65240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12131 n_87400_65240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12132 n_92340_76440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12133 n_88920_87640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12134 n_85880_87640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12135 n_83600_51240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12136 n_85500_51240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12137 n_90820_56840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12138 n_92720_59640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12139 n_90820_82040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12140 n_77900_87640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12141 n_82080_54040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12142 n_80560_56840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12143 n_82080_56840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12144 n_78660_56840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12145 n_76380_54040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12146 n_76760_65240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12147 n_76760_56840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12148 n_78660_65240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12149 n_77900_68040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12150 n_79040_68040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12151 n_62320_82040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12152 n_70300_87640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12153 n_73720_82040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12154 n_72200_84840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12155 n_82080_51240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12156 n_86260_54040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12157 n_87400_48440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12158 n_85500_59640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12159 n_80560_68040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12160 n_77140_70840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12161 n_80560_70840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12162 n_80560_73640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12163 n_78660_79240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12164 n_78280_82040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12165 n_80180_82040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12166 n_76760_84840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12167 n_78660_84840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12168 n_67260_51240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12169 n_70300_51240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12170 n_68020_54040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12171 n_49780_54040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12172 n_50920_51240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12173 n_52060_51240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12174 n_66120_51240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12175 n_79040_51240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12176 n_87400_51240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12177 n_49400_48440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12178 n_51680_45640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12179 n_53200_48440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12180 n_65360_42840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12181 n_70300_42840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12182 n_92720_42840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12183 n_50540_42840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12184 n_45220_42840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12185 n_46740_45640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12186 n_61560_40040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12187 n_85500_42840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12188 n_42940_48440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12189 n_53200_45640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12190 n_73720_45640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12191 n_73340_40040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12192 n_53200_42840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12193 n_44080_48440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12194 n_49780_56840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12195 n_48260_62440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12196 n_52060_54040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12197 n_48260_65240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12198 n_49780_62440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12199 n_59660_62440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12200 n_44840_73640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12201 n_50920_68040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12202 n_72200_56840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12203 n_56620_65240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12204 n_61560_62440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12205 n_58520_65240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12206 n_60420_65240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12207 n_73720_62440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12208 n_63460_68040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12209 n_76380_62440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12210 n_63080_82040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12211 n_75240_59640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12212 n_77520_62440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12213 n_73340_59640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12214 n_69160_62440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12215 n_49400_73640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12216 n_55860_68040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12217 n_46740_73640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12218 n_46360_76440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12219 n_40660_76440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12220 n_48260_73640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12221 n_40660_70840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12222 n_49780_76440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12223 n_50920_79240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12224 n_58520_68040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12225 n_61560_73640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12226 n_66880_73640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12227 n_74100_68040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12228 n_75240_68040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12229 n_72960_68040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12230 n_68020_62440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12231 n_55480_48440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12232 n_68780_70840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12233 n_48260_76440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12234 n_47500_79240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12235 n_48640_79240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12236 n_58520_70840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12237 n_60040_76440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12238 n_60420_70840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12239 n_63080_73640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12240 n_71820_73640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12241 n_76760_73640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12242 n_60040_79240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12243 n_63080_79240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12244 n_67260_70840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12245 n_58140_51240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12246 n_70300_48440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12247 n_40660_79240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12248 n_40280_82040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12249 n_43700_79240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12250 n_40280_87640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12251 n_63080_76440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12252 n_50920_82040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12253 n_53580_82040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12254 n_65740_73640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12255 n_70300_76440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12256 n_40280_84840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12257 n_41420_87640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12258 n_46740_87640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12259 n_46740_84840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12260 n_61940_84840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12261 n_63080_84840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12262 n_49400_84840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12263 n_55100_82040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12264 n_46740_51240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12265 n_43320_68040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12266 n_43320_76440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12267 n_44080_82040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12268 n_65360_62440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12269 n_66880_62440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12270 n_65360_56840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12271 n_63080_54040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12272 n_68780_56840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12273 n_67260_82040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12274 n_65740_82040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12275 n_58520_84840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12276 n_64600_84840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12277 n_65360_65240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12278 n_67260_65240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12279 n_63460_59640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12280 n_63460_56840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12281 n_60040_54040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12282 n_68780_59640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12283 n_66880_59640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12284 n_70300_59640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12285 n_70300_56840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12286 n_70300_65240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12287 n_68400_65240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12288 n_71820_65240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12289 n_71820_68040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12290 n_70300_68040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12291 n_71820_70840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12292 n_68780_76440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12293 n_55100_79240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12294 n_59660_82040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12295 n_56240_82040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12296 n_87400_62440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12297 n_87020_59640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12298 n_85880_62440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12299 n_83220_65240 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12300 n_84740_62440 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12301 n_83220_68040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12302 n_83600_70840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12303 n_83220_73640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12304 n_85500_82040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12305 n_71060_82040 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12306 n_44460_56840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12307 n_60040_56840 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12308 n_60040_59640 0 PWL(106000ps 0uA 106030ps 0uA 106031ps 30uA 106059ps 30uA 106060ps 0uA)
I12309 n_90820_68040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12310 n_91200_70840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12311 n_93480_79240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12312 n_91960_87640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12313 n_90440_62440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12314 n_93480_68040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12315 n_93480_73640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12316 n_93480_76440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12317 n_54720_48440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12318 n_56240_48440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12319 n_61940_48440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12320 n_40660_56840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12321 n_79040_42840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12322 n_93480_48440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12323 n_92340_48440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12324 n_50920_48440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12325 n_70300_40040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12326 n_91580_40040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12327 n_87020_40040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12328 n_88160_40040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12329 n_52440_40040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12330 n_90440_40040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12331 n_40280_40040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12332 n_60040_45640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12333 n_79040_40040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12334 n_77140_40040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12335 n_55100_40040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12336 n_40660_51240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12337 n_44460_68040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12338 n_45600_68040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12339 n_43320_62440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12340 n_44460_62440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12341 n_47500_68040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12342 n_46740_65240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12343 n_44840_51240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12344 n_54720_42840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12345 n_74860_40040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12346 n_76760_42840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12347 n_56620_45640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12348 n_41420_40040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12349 n_83600_42840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12350 n_51680_42840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12351 n_83600_40040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12352 n_87020_45640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12353 n_92720_40040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12354 n_68400_40040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12355 n_51680_48440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12356 n_85120_48440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12357 n_90440_48440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12358 n_78280_48440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12359 n_41420_54040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12360 n_60040_48440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12361 n_55100_54040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12362 n_54720_51240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12363 n_90440_76440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12364 n_90440_73640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12365 n_92340_65240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12366 n_90820_59640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12367 n_87400_84840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12368 n_91580_79240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12369 n_87400_73640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12370 n_88540_68040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12371 n_83220_54040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12372 n_91200_54040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12373 n_92340_56840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12374 n_90820_65240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12375 n_87400_65240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12376 n_87400_76440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12377 n_92340_76440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12378 n_88920_82040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12379 n_88920_87640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12380 n_85880_87640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12381 n_83600_51240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12382 n_85500_51240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12383 n_77520_54040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12384 n_87400_79240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12385 n_92720_59640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12386 n_88920_65240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12387 n_92340_73640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12388 n_88920_76440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12389 n_79040_54040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12390 n_80560_54040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12391 n_82080_54040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12392 n_76760_56840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12393 n_78280_70840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12394 n_70300_79240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12395 n_67260_84840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12396 n_88920_79240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12397 n_67260_87640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12398 n_65360_87640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12399 n_68780_87640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12400 n_71820_87640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12401 n_70300_87640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12402 n_72200_84840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12403 n_82080_51240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12404 n_87400_48440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12405 n_85500_59640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12406 n_80560_68040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12407 n_77140_70840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12408 n_76760_76440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12409 n_72200_76440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12410 n_76760_79240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12411 n_80560_79240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12412 n_70300_51240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12413 n_68020_54040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12414 n_61940_51240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12415 n_52060_51240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12416 n_79040_51240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12417 n_87400_51240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12418 n_83600_48440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12419 n_53200_48440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12420 n_70300_42840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12421 n_92720_42840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12422 n_90440_45640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12423 n_85500_40040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12424 n_50540_42840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12425 n_85500_42840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12426 n_43320_40040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12427 n_53200_45640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12428 n_76760_45640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12429 n_73340_40040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12430 n_53200_42840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12431 n_43320_51240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12432 n_57000_54040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12433 n_52060_54040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12434 n_61560_65240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12435 n_58520_65240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12436 n_59660_68040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12437 n_60420_65240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12438 n_73720_62440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12439 n_66880_68040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12440 n_63460_68040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12441 n_63080_65240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12442 n_75240_62440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12443 n_76380_59640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12444 n_61940_68040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12445 n_55100_56840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12446 n_69160_62440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12447 n_50920_73640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12448 n_49400_73640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12449 n_46740_73640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12450 n_46360_76440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12451 n_40660_76440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12452 n_40660_70840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12453 n_61560_73640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12454 n_66880_73640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12455 n_63460_70840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12456 n_74100_68040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12457 n_65360_68040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12458 n_68780_68040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12459 n_75240_65240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12460 n_68020_62440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12461 n_68780_70840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12462 n_53580_65240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12463 n_53580_68040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12464 n_54720_68040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12465 n_48260_76440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12466 n_47500_79240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12467 n_48640_79240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12468 n_58520_70840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12469 n_60040_76440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12470 n_60420_70840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12471 n_63080_73640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12472 n_60040_79240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12473 n_63080_79240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12474 n_67260_70840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12475 n_58140_51240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12476 n_46360_68040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12477 n_44840_70840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12478 n_44840_76440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12479 n_40660_79240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12480 n_40280_82040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12481 n_43700_79240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12482 n_40280_87640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12483 n_63080_76440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12484 n_50920_82040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12485 n_53580_82040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12486 n_52820_79240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12487 n_44080_59640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12488 n_42940_82040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12489 n_45220_82040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12490 n_40280_84840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12491 n_41420_87640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12492 n_46740_87640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12493 n_46740_84840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12494 n_49400_84840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12495 n_55100_82040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12496 n_42940_54040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12497 n_73340_87640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12498 n_70300_65240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12499 n_68400_65240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12500 n_71820_65240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12501 n_71820_68040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12502 n_70300_68040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12503 n_71820_70840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12504 n_68780_76440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12505 n_55100_79240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12506 n_88160_59640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12507 n_84740_62440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12508 n_85500_70840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12509 n_84740_73640 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12510 n_85880_68040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12511 n_83600_76440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12512 n_85500_76440 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12513 n_85500_79240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12514 n_83600_82040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12515 n_83600_79240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12516 n_85500_82040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12517 n_69920_82040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12518 n_68780_82040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12519 n_71060_82040 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12520 n_43320_65240 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12521 n_44460_56840 0 PWL(108000ps 0uA 108030ps 0uA 108031ps 30uA 108059ps 30uA 108060ps 0uA)
I12522 n_93480_62440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12523 n_93480_79240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12524 n_93100_87640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12525 n_90440_62440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12526 n_93480_68040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12527 n_93100_84840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12528 n_84740_87640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12529 n_65740_45640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12530 n_61940_48440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12531 n_40280_54040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12532 n_93480_54040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12533 n_92340_48440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12534 n_41800_42840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12535 n_70300_40040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12536 n_87020_40040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12537 n_88160_40040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12538 n_52440_40040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12539 n_40660_42840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12540 n_56620_40040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12541 n_93480_45640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12542 n_40280_48440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12543 n_60040_45640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12544 n_72200_40040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12545 n_40660_51240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12546 n_44460_68040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12547 n_45600_68040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12548 n_47500_68040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12549 n_46740_65240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12550 n_44840_51240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12551 n_71820_42840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12552 n_56620_45640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12553 n_41420_48440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12554 n_88920_45640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12555 n_57760_40040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12556 n_43700_42840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12557 n_51680_42840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12558 n_83600_40040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12559 n_87020_45640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12560 n_68400_40040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12561 n_48260_45640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12562 n_85120_48440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12563 n_92340_51240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12564 n_47880_54040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12565 n_60040_48440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12566 n_64600_51240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12567 n_81700_87640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12568 n_90820_84840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12569 n_92340_65240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12570 n_90820_59640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12571 n_90060_87640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12572 n_91580_79240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12573 n_91580_62440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12574 n_83220_54040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12575 n_91200_54040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12576 n_90820_65240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12577 n_88920_70840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12578 n_87400_65240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12579 n_87400_70840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12580 n_87400_76440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12581 n_92340_76440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12582 n_87780_87640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12583 n_88920_82040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12584 n_85880_87640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12585 n_83600_51240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12586 n_80560_51240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12587 n_84740_54040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12588 n_77520_54040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12589 n_87400_79240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12590 n_92720_59640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12591 n_88920_65240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12592 n_88920_76440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12593 n_90060_79240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12594 n_90820_82040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12595 n_79040_87640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12596 n_79040_54040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12597 n_80560_54040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12598 n_82080_54040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12599 n_80560_65240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12600 n_77900_68040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12601 n_76000_70840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12602 n_79040_68040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12603 n_78280_70840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12604 n_74860_70840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12605 n_73720_70840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12606 n_75240_76440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12607 n_73720_73640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12608 n_62320_82040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12609 n_65360_87640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12610 n_72200_84840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12611 n_85500_56840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12612 n_82080_59640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12613 n_85500_59640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12614 n_84740_65240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12615 n_82080_65240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12616 n_82080_68040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12617 n_82080_70840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12618 n_81700_73640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12619 n_80560_70840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12620 n_78660_73640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12621 n_78660_76440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12622 n_78660_79240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12623 n_72200_76440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12624 n_78280_82040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12625 n_76760_79240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12626 n_80560_79240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12627 n_76760_84840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12628 n_78660_84840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12629 n_74860_84840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12630 n_68780_51240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12631 n_61940_51240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12632 n_49780_54040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12633 n_90820_51240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12634 n_83600_48440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12635 n_49400_48440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12636 n_70300_42840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12637 n_90440_45640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12638 n_85500_40040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12639 n_50540_42840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12640 n_45220_42840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12641 n_61560_40040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12642 n_88920_42840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12643 n_42940_48440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12644 n_53200_45640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12645 n_73720_45640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12646 n_43320_51240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12647 n_57000_54040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12648 n_52060_54040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12649 n_66880_68040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12650 n_60800_68040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12651 n_60040_73640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12652 n_77520_62440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12653 n_59660_70840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12654 n_55100_56840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12655 n_69160_62440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12656 n_50920_73640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12657 n_49400_73640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12658 n_46740_73640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12659 n_46360_76440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12660 n_40660_76440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12661 n_40660_70840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12662 n_58520_68040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12663 n_58520_73640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12664 n_70300_73640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12665 n_63460_70840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12666 n_65360_68040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12667 n_68780_68040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12668 n_68020_62440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12669 n_55480_48440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12670 n_53580_65240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12671 n_53580_68040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12672 n_54720_68040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12673 n_48260_76440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12674 n_47500_79240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12675 n_48640_79240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12676 n_58520_70840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12677 n_60040_76440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12678 n_60420_70840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12679 n_71820_73640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12680 n_60040_79240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12681 n_63080_79240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12682 n_58140_51240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12683 n_46360_68040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12684 n_44840_70840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12685 n_44840_76440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12686 n_41800_70840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12687 n_43700_79240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12688 n_63080_76440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12689 n_80560_76440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12690 n_50920_82040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12691 n_49400_82040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12692 n_54720_84840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12693 n_53580_82040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12694 n_47500_56840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12695 n_52820_79240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12696 n_46740_84840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12697 n_61940_84840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12698 n_49400_84840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12699 n_55100_82040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12700 n_73340_87640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12701 n_71820_68040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12702 n_73720_65240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12703 n_70300_68040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12704 n_68780_76440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12705 n_88160_59640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12706 n_85880_62440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12707 n_83220_65240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12708 n_83220_62440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12709 n_83220_68040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12710 n_83600_70840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12711 n_85500_70840 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12712 n_83220_73640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12713 n_84740_73640 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12714 n_85880_68040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12715 n_83600_76440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12716 n_85500_76440 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12717 n_85500_79240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12718 n_83600_82040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12719 n_83600_79240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12720 n_69920_82040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12721 n_68780_82040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12722 n_71060_82040 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12723 n_43320_65240 0 PWL(110000ps 0uA 110030ps 0uA 110031ps 30uA 110059ps 30uA 110060ps 0uA)
I12724 n_93480_79240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12725 n_93100_87640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12726 n_93480_56840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12727 n_90440_62440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12728 n_93480_68040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12729 n_93100_84840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12730 n_83600_87640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12731 n_61940_48440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12732 n_40660_56840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12733 n_92340_48440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12734 n_50920_48440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12735 n_63840_40040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12736 n_70300_40040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12737 n_87020_40040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12738 n_88160_40040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12739 n_42940_42840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12740 n_93480_45640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12741 n_80560_40040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12742 n_46360_40040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12743 n_40280_40040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12744 n_40280_48440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12745 n_60040_45640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12746 n_79040_40040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12747 n_77140_40040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12748 n_40660_51240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12749 n_44840_51240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12750 n_74860_40040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12751 n_76760_42840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12752 n_56620_45640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12753 n_41420_48440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12754 n_41420_40040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12755 n_49400_40040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12756 n_80180_42840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12757 n_88920_45640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12758 n_44840_45640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12759 n_83600_40040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12760 n_87020_45640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12761 n_68400_40040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12762 n_63460_42840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12763 n_51680_48440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12764 n_85120_48440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12765 n_41420_54040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12766 n_60040_48440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12767 n_80180_87640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12768 n_90820_84840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12769 n_92340_65240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12770 n_90820_59640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12771 n_88920_56840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12772 n_90060_87640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12773 n_91580_79240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12774 n_92720_82040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12775 n_88920_87640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12776 n_80560_51240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12777 n_85500_51240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12778 n_84740_54040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12779 n_90820_56840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12780 n_92720_59640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12781 n_91960_68040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12782 n_90820_82040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12783 n_77900_87640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12784 n_80560_56840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12785 n_82080_56840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12786 n_78660_56840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12787 n_83600_56840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12788 n_76760_65240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12789 n_78660_65240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12790 n_80560_65240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12791 n_79040_68040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12792 n_78280_70840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12793 n_75240_73640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12794 n_75240_76440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12795 n_73720_79240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12796 n_70300_79240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12797 n_67260_84840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12798 n_65740_84840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12799 n_65360_87640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12800 n_68780_87640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12801 n_71820_87640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12802 n_70300_87640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12803 n_72200_84840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12804 n_82080_51240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12805 n_85500_56840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12806 n_87400_48440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12807 n_82080_59640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12808 n_82080_65240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12809 n_81700_76440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12810 n_72200_76440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12811 n_74860_84840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12812 n_61940_51240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12813 n_52060_51240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12814 n_83600_48440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12815 n_53200_48440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12816 n_65360_42840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12817 n_70300_42840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12818 n_90440_45640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12819 n_85500_40040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12820 n_46740_45640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12821 n_88920_42840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12822 n_82080_42840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12823 n_51300_40040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12824 n_43320_40040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12825 n_42940_48440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12826 n_53200_45640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12827 n_76760_45640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12828 n_73340_40040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12829 n_43320_51240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12830 n_52060_54040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12831 n_77520_62440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12832 n_66880_73640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12833 n_58140_79240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12834 n_55480_48440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12835 n_68780_70840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12836 n_56620_79240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12837 n_60040_79240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12838 n_63080_79240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12839 n_65740_76440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12840 n_67260_70840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12841 n_70300_48440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12842 n_57380_76440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12843 n_63080_76440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12844 n_65740_73640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12845 n_73340_87640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12846 n_71820_68040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12847 n_73720_65240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12848 n_70300_70840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12849 n_67260_76440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12850 n_68780_76440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12851 n_65740_79240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12852 n_64600_79240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12853 n_64600_76440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12854 n_87400_62440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12855 n_87020_59640 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12856 n_85880_62440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12857 n_83220_65240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12858 n_83220_62440 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12859 n_83220_68040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12860 n_83600_70840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12861 n_85500_70840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12862 n_85880_68040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12863 n_85500_82040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12864 n_69920_82040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12865 n_68780_82040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12866 n_71060_82040 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12867 n_43320_65240 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12868 n_44460_56840 0 PWL(112000ps 0uA 112030ps 0uA 112031ps 30uA 112059ps 30uA 112060ps 0uA)
I12869 n_91200_70840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12870 n_93480_79240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12871 n_93480_68040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12872 n_93480_76440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12873 n_83600_87640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12874 n_84740_87640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12875 n_65740_45640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12876 n_61940_48440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12877 n_93480_54040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12878 n_92340_48440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12879 n_40660_42840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12880 n_42940_42840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12881 n_90440_40040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12882 n_40280_40040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12883 n_82080_48440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12884 n_55100_40040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12885 n_40660_51240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12886 n_50160_59640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12887 n_42180_73640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12888 n_44460_68040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12889 n_45600_68040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12890 n_40660_65240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12891 n_41800_68040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12892 n_47500_68040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12893 n_46740_65240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12894 n_52060_73640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12895 n_51300_59640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12896 n_44840_51240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12897 n_54720_42840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12898 n_80180_45640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12899 n_41420_40040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12900 n_83600_42840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12901 n_44840_45640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12902 n_43700_42840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12903 n_85120_48440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12904 n_92340_51240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12905 n_60040_48440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12906 n_64600_51240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12907 n_81700_87640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12908 n_80180_87640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12909 n_90440_76440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12910 n_92340_65240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12911 n_91580_79240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12912 n_87400_73640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12913 n_87400_70840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12914 n_92720_82040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12915 n_80560_51240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12916 n_85500_51240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12917 n_84740_54040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12918 n_91960_68040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12919 n_90060_79240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12920 n_77900_87640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12921 n_79040_87640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12922 n_79040_68040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12923 n_78280_70840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12924 n_74860_70840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12925 n_73720_70840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12926 n_88920_79240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12927 n_67260_87640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12928 n_65360_87640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12929 n_72200_84840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12930 n_82080_51240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12931 n_85500_56840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12932 n_87400_48440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12933 n_82080_59640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12934 n_82080_65240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12935 n_85880_65240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12936 n_87400_68040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12937 n_80560_73640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12938 n_81700_76440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12939 n_72200_76440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12940 n_74860_82040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12941 n_76760_82040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12942 n_68780_51240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12943 n_61940_51240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12944 n_90820_51240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12945 n_83600_48440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12946 n_45220_42840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12947 n_46740_45640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12948 n_85500_42840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12949 n_43320_40040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12950 n_82080_45640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12951 n_53200_42840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12952 n_43320_51240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12953 n_57000_54040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12954 n_52060_54040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12955 n_48260_65240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12956 n_59660_62440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12957 n_50920_68040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12958 n_53580_59640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12959 n_53580_62440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12960 n_52060_65240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12961 n_49400_65240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12962 n_56620_65240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12963 n_61560_62440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12964 n_61560_65240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12965 n_59660_68040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12966 n_60800_68040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12967 n_60040_73640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12968 n_63080_65240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12969 n_77520_62440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12970 n_61940_68040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12971 n_59660_70840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12972 n_55100_56840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12973 n_55100_70840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12974 n_53580_70840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12975 n_50920_70840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12976 n_50920_73640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12977 n_49400_73640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12978 n_55860_68040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12979 n_46360_76440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12980 n_48260_73640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12981 n_49780_76440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12982 n_50920_79240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12983 n_58520_73640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12984 n_70300_73640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12985 n_66880_73640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12986 n_58140_79240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12987 n_68780_70840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12988 n_53580_65240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12989 n_53580_68040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12990 n_49400_70840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12991 n_46740_70840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12992 n_48260_76440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12993 n_47500_79240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12994 n_48640_79240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12995 n_58520_70840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12996 n_60040_76440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12997 n_60420_70840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12998 n_71820_73640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I12999 n_60040_79240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13000 n_63080_79240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13001 n_52060_82040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13002 n_65740_76440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13003 n_67260_70840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13004 n_58140_51240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13005 n_70300_48440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13006 n_46360_68040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13007 n_44840_70840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13008 n_43320_70840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13009 n_40280_82040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13010 n_43700_79240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13011 n_40280_87640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13012 n_63080_76440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13013 n_50920_82040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13014 n_53580_82040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13015 n_65740_73640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13016 n_52820_79240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13017 n_45220_82040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13018 n_42940_84840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13019 n_40280_84840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13020 n_41420_87640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13021 n_46740_87640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13022 n_46740_84840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13023 n_49400_84840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13024 n_55100_82040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13025 n_42940_54040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13026 n_43320_68040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13027 n_43320_76440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13028 n_44080_82040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13029 n_65360_62440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13030 n_65360_54040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13031 n_65360_56840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13032 n_68780_56840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13033 n_73340_87640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13034 n_65360_65240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13035 n_63460_62440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13036 n_63460_59640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13037 n_63460_56840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13038 n_68780_59640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13039 n_70300_59640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13040 n_70300_56840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13041 n_71820_59640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13042 n_70300_65240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13043 n_71820_65240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13044 n_71820_68040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13045 n_70300_70840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13046 n_67260_76440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13047 n_68780_76440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13048 n_64600_79240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13049 n_53960_79240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13050 n_64600_76440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13051 n_85880_62440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13052 n_83220_65240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13053 n_83220_62440 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13054 n_83220_68040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13055 n_84740_68040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13056 n_83600_70840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13057 n_85500_70840 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13058 n_85880_68040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13059 n_85880_73640 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13060 n_81700_79240 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13061 n_69920_82040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13062 n_71060_82040 0 PWL(114000ps 0uA 114030ps 0uA 114031ps 30uA 114059ps 30uA 114060ps 0uA)
I13063 n_93480_79240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13064 n_91960_87640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13065 n_90440_62440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13066 n_93480_68040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13067 n_61940_48440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13068 n_40280_54040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13069 n_92340_48440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13070 n_41800_42840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13071 n_91580_40040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13072 n_88160_40040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13073 n_40660_42840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13074 n_56620_40040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13075 n_90440_40040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13076 n_46360_40040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13077 n_40280_40040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13078 n_60040_45640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13079 n_82080_48440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13080 n_77140_40040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13081 n_40660_51240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13082 n_43320_59640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13083 n_50160_59640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13084 n_42180_73640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13085 n_44460_68040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13086 n_45600_68040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13087 n_43320_62440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13088 n_44460_62440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13089 n_47500_68040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13090 n_46740_65240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13091 n_52060_73640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13092 n_51300_59640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13093 n_46740_59640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13094 n_44840_51240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13095 n_74860_40040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13096 n_80180_45640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13097 n_56620_45640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13098 n_41420_40040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13099 n_49400_40040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13100 n_83600_42840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13101 n_57760_40040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13102 n_43700_42840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13103 n_83600_40040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13104 n_92720_40040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13105 n_48260_45640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13106 n_85120_48440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13107 n_47880_54040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13108 n_60040_48440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13109 n_92340_65240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13110 n_90820_59640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13111 n_87400_84840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13112 n_91580_79240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13113 n_92720_82040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13114 n_87780_87640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13115 n_80560_51240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13116 n_85500_51240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13117 n_84740_54040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13118 n_92720_59640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13119 n_91960_68040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13120 n_78660_56840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13121 n_76760_65240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13122 n_78660_65240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13123 n_80560_65240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13124 n_79040_68040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13125 n_78280_70840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13126 n_71820_79240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13127 n_65740_84840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13128 n_62320_82040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13129 n_82080_51240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13130 n_85500_56840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13131 n_87400_48440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13132 n_85500_59640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13133 n_84740_65240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13134 n_82080_68040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13135 n_85880_65240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13136 n_87400_68040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13137 n_82080_70840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13138 n_80560_70840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13139 n_80560_73640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13140 n_81700_76440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13141 n_78660_73640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13142 n_78660_76440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13143 n_78660_79240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13144 n_72200_76440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13145 n_78280_82040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13146 n_76760_84840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13147 n_78660_84840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13148 n_61940_51240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13149 n_49780_54040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13150 n_83600_48440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13151 n_49400_48440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13152 n_92720_42840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13153 n_85500_40040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13154 n_45220_42840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13155 n_61560_40040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13156 n_85500_42840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13157 n_51300_40040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13158 n_43320_40040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13159 n_53200_45640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13160 n_82080_45640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13161 n_73340_40040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13162 n_43320_51240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13163 n_57000_54040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13164 n_49780_56840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13165 n_48260_62440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13166 n_52060_54040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13167 n_49780_62440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13168 n_44840_73640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13169 n_53580_59640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13170 n_53580_62440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13171 n_52060_65240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13172 n_49400_65240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13173 n_55100_56840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13174 n_55100_70840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13175 n_53580_70840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13176 n_50920_70840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13177 n_50920_73640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13178 n_46740_73640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13179 n_40660_76440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13180 n_40660_70840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13181 n_55480_48440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13182 n_53580_65240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13183 n_53580_68040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13184 n_49400_70840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13185 n_46740_70840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13186 n_56620_79240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13187 n_60040_79240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13188 n_63080_79240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13189 n_52060_82040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13190 n_46360_68040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13191 n_44840_70840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13192 n_43320_70840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13193 n_41800_70840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13194 n_40280_82040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13195 n_40280_87640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13196 n_57380_76440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13197 n_63080_76440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13198 n_49400_82040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13199 n_54720_84840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13200 n_44080_59640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13201 n_42940_82040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13202 n_42940_84840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13203 n_40280_84840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13204 n_41420_87640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13205 n_46740_87640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13206 n_61940_84840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13207 n_68780_76440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13208 n_65740_79240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13209 n_53960_79240 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13210 n_85880_62440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13211 n_84740_62440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13212 n_83220_62440 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13213 n_83220_68040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13214 n_84740_68040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13215 n_83600_70840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13216 n_85500_70840 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13217 n_85880_68040 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13218 n_85880_73640 0 PWL(116000ps 0uA 116030ps 0uA 116031ps 30uA 116059ps 30uA 116060ps 0uA)
I13219 n_87020_87640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13220 n_93100_87640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13221 n_93480_68040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13222 n_93480_76440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13223 n_93100_84840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13224 n_44080_54040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13225 n_40660_56840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13226 n_48640_40040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13227 n_50920_48440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13228 n_52440_40040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13229 n_40660_42840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13230 n_42940_42840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13231 n_56620_40040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13232 n_93480_45640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13233 n_72200_40040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13234 n_40660_45640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13235 n_40660_51240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13236 n_43320_59640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13237 n_46740_59640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13238 n_44840_51240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13239 n_45220_48440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13240 n_71820_42840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13241 n_88920_45640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13242 n_57760_40040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13243 n_44840_45640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13244 n_43700_42840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13245 n_51680_42840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13246 n_51680_48440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13247 n_47880_42840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13248 n_41420_54040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13249 n_49020_51240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13250 n_90820_84840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13251 n_90440_76440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13252 n_92340_65240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13253 n_90060_87640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13254 n_85120_84840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13255 n_83600_84840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13256 n_88920_87640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13257 n_80560_51240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13258 n_84740_54040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13259 n_91960_68040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13260 n_90060_79240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13261 n_90820_82040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13262 n_76000_70840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13263 n_79040_68040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13264 n_78280_70840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13265 n_75240_73640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13266 n_73720_79240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13267 n_70300_79240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13268 n_67260_84840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13269 n_71820_79240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13270 n_88920_79240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13271 n_67260_87640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13272 n_68780_87640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13273 n_68780_84840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13274 n_70300_84840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13275 n_73720_82040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13276 n_85500_56840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13277 n_85500_59640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13278 n_84740_65240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13279 n_82080_68040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13280 n_85880_65240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13281 n_87400_68040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13282 n_82080_70840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13283 n_80560_70840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13284 n_80560_73640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13285 n_81700_76440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13286 n_78660_73640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13287 n_78660_76440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13288 n_78660_79240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13289 n_78280_82040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13290 n_80180_82040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13291 n_74860_82040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13292 n_76760_82040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13293 n_50920_51240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13294 n_52060_51240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13295 n_51680_45640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13296 n_53200_48440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13297 n_50540_42840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13298 n_45220_42840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13299 n_46740_45640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13300 n_61560_40040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13301 n_88920_42840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13302 n_73720_45640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13303 n_44080_48440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13304 n_43320_51240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13305 n_57000_54040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13306 n_49780_56840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13307 n_48260_62440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13308 n_48260_65240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13309 n_49780_62440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13310 n_59660_62440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13311 n_44840_73640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13312 n_50920_68040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13313 n_56620_65240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13314 n_61560_62440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13315 n_61560_65240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13316 n_59660_68040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13317 n_60800_68040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13318 n_60040_73640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13319 n_63080_65240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13320 n_61940_68040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13321 n_59660_70840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13322 n_49400_73640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13323 n_55860_68040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13324 n_46740_73640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13325 n_46360_76440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13326 n_40660_76440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13327 n_48260_73640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13328 n_40660_70840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13329 n_49780_76440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13330 n_50920_79240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13331 n_58520_73640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13332 n_56620_73640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13333 n_58140_79240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13334 n_55480_48440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13335 n_48260_76440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13336 n_47500_79240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13337 n_48640_79240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13338 n_58520_70840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13339 n_60040_76440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13340 n_60420_70840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13341 n_63080_73640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13342 n_56620_79240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13343 n_52060_82040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13344 n_40660_79240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13345 n_40280_82040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13346 n_43700_79240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13347 n_44080_84840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13348 n_40280_87640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13349 n_57380_76440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13350 n_80560_76440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13351 n_49400_82040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13352 n_47120_82040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13353 n_50160_84840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13354 n_41420_87640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13355 n_46740_87640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13356 n_46740_84840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13357 n_49400_87640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13358 n_64220_82040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13359 n_65360_62440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13360 n_65360_54040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13361 n_65360_56840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13362 n_68780_56840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13363 n_45220_87640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13364 n_51680_84840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13365 n_67260_82040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13366 n_65360_65240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13367 n_63460_62440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13368 n_63460_59640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13369 n_63460_56840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13370 n_68780_59640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13371 n_70300_59640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13372 n_70300_56840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13373 n_71820_59640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13374 n_70300_65240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13375 n_71820_65240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13376 n_71820_68040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13377 n_70300_70840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13378 n_67260_76440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13379 n_65740_79240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13380 n_64600_79240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13381 n_57380_82040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13382 n_58520_82040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13383 n_59660_82040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13384 n_88920_62440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13385 n_85880_62440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13386 n_84740_62440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13387 n_83220_62440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13388 n_83220_68040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13389 n_84740_68040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13390 n_83600_70840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13391 n_85500_70840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13392 n_85880_68040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13393 n_85880_73640 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13394 n_83600_76440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13395 n_81700_79240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13396 n_85500_76440 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13397 n_85500_79240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13398 n_83600_79240 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13399 n_85500_82040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13400 n_68780_82040 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13401 n_44460_56840 0 PWL(118000ps 0uA 118030ps 0uA 118031ps 30uA 118059ps 30uA 118060ps 0uA)
I13402 n_92340_54040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13403 n_93480_62440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13404 n_91200_70840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13405 n_93100_87640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13406 n_93480_56840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13407 n_90440_62440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13408 n_93480_73640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13409 n_93480_76440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13410 n_93100_84840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13411 n_65740_40040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13412 n_54720_48440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13413 n_56240_48440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13414 n_44080_54040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13415 n_40660_56840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13416 n_79040_42840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13417 n_93480_48440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13418 n_41800_42840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13419 n_48640_40040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13420 n_50920_48440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13421 n_63840_40040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13422 n_70300_40040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13423 n_91580_40040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13424 n_87020_40040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13425 n_52440_40040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13426 n_42940_42840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13427 n_56620_40040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13428 n_90440_40040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13429 n_77140_40040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13430 n_40660_45640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13431 n_43320_59640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13432 n_42180_73640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13433 n_40660_65240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13434 n_47500_40040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13435 n_89300_48440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13436 n_41800_68040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13437 n_52060_73640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13438 n_46740_59640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13439 n_45220_48440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13440 n_74860_40040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13441 n_83600_42840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13442 n_57760_40040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13443 n_44840_45640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13444 n_51680_42840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13445 n_87020_45640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13446 n_92720_40040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13447 n_68400_40040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13448 n_63460_42840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13449 n_51680_48440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13450 n_47880_42840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13451 n_48260_45640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13452 n_90440_48440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13453 n_78280_48440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13454 n_41420_54040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13455 n_49020_51240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13456 n_55100_54040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13457 n_54720_51240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13458 n_63080_51240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13459 n_90820_84840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13460 n_90440_76440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13461 n_90440_73640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13462 n_90820_59640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13463 n_88920_56840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13464 n_90060_87640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13465 n_87400_73640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13466 n_91580_62440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13467 n_89300_54040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13468 n_73340_51240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13469 n_71820_48440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13470 n_73340_48440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13471 n_73720_54040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13472 n_88920_51240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13473 n_83220_54040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13474 n_91200_54040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13475 n_90820_65240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13476 n_88920_70840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13477 n_87400_65240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13478 n_87400_76440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13479 n_92720_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13480 n_92340_76440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13481 n_83600_84840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13482 n_82080_84840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13483 n_85880_87640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13484 n_83600_51240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13485 n_80560_51240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13486 n_85500_51240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13487 n_84740_54040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13488 n_90820_56840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13489 n_92720_59640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13490 n_92340_73640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13491 n_90060_79240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13492 n_90820_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13493 n_79040_54040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13494 n_80560_54040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13495 n_82080_54040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13496 n_80560_56840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13497 n_80180_59640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13498 n_78660_56840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13499 n_83600_56840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13500 n_76380_54040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13501 n_76760_65240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13502 n_78660_65240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13503 n_80560_65240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13504 n_76000_70840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13505 n_79040_68040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13506 n_75240_73640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13507 n_73720_70840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13508 n_73720_79240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13509 n_70300_79240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13510 n_67260_84840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13511 n_88920_79240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13512 n_67260_87640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13513 n_68780_87640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13514 n_68780_84840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13515 n_70300_87640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13516 n_70300_84840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13517 n_73720_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13518 n_82080_51240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13519 n_85500_56840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13520 n_82080_59640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13521 n_85500_59640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13522 n_84740_65240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13523 n_82080_65240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13524 n_82080_68040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13525 n_85880_65240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13526 n_87400_68040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13527 n_82080_70840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13528 n_80560_68040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13529 n_77140_70840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13530 n_81700_73640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13531 n_80560_73640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13532 n_78660_73640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13533 n_78660_76440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13534 n_78660_79240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13535 n_76760_76440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13536 n_72200_76440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13537 n_78280_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13538 n_80180_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13539 n_74860_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13540 n_76760_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13541 n_60800_51240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13542 n_71820_51240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13543 n_71820_54040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13544 n_53200_51240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13545 n_68020_54040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13546 n_59280_51240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13547 n_61940_51240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13548 n_50920_51240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13549 n_41800_56840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13550 n_75240_54040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13551 n_76380_51240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13552 n_76760_48440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13553 n_87400_51240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13554 n_83600_48440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13555 n_85500_45640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13556 n_50160_45640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13557 n_51680_45640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13558 n_48260_48440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13559 n_61560_42840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13560 n_70300_42840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13561 n_89300_40040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13562 n_90440_45640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13563 n_85500_40040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13564 n_81700_40040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13565 n_50540_42840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13566 n_46740_45640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13567 n_61560_40040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13568 n_68020_48440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13569 n_68780_45640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13570 n_85500_42840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13571 n_82080_42840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13572 n_73720_42840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13573 n_53200_45640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13574 n_58520_45640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13575 n_82080_45640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13576 n_80560_48440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13577 n_73340_40040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13578 n_44080_48440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13579 n_57000_54040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13580 n_48640_59640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13581 n_52060_54040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13582 n_40280_59640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13583 n_72200_56840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13584 n_61560_62440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13585 n_61560_65240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13586 n_58520_65240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13587 n_59660_68040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13588 n_60420_65240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13589 n_73720_62440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13590 n_60800_68040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13591 n_63460_68040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13592 n_63080_65240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13593 n_75240_62440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13594 n_76380_59640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13595 n_75240_59640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13596 n_72200_62440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13597 n_53580_73640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13598 n_50920_73640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13599 n_49400_73640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13600 n_55860_68040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13601 n_46740_73640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13602 n_46360_76440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13603 n_40660_76440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13604 n_40660_70840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13605 n_46360_79240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13606 n_58520_68040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13607 n_70300_73640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13608 n_56620_73640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13609 n_58140_79240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13610 n_74100_68040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13611 n_75240_65240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13612 n_40280_73640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13613 n_45600_84840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13614 n_49400_79240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13615 n_63080_73640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13616 n_71820_73640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13617 n_56620_79240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13618 n_60040_79240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13619 n_63080_79240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13620 n_52060_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13621 n_58140_51240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13622 n_40660_79240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13623 n_40280_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13624 n_43700_79240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13625 n_44080_84840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13626 n_40280_87640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13627 n_57380_76440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13628 n_63080_76440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13629 n_50920_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13630 n_49400_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13631 n_47120_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13632 n_53580_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13633 n_50160_84840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13634 n_52820_79240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13635 n_43320_87640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13636 n_49400_84840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13637 n_52440_87640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13638 n_49400_87640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13639 n_64220_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13640 n_58140_87640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13641 n_55100_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13642 n_42940_54040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13643 n_46740_51240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13644 n_41800_65240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13645 n_65360_59640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13646 n_65360_62440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13647 n_65360_54040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13648 n_65360_56840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13649 n_68780_56840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13650 n_59280_87640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13651 n_60800_84840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13652 n_61180_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13653 n_54340_76440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13654 n_54340_87640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13655 n_67260_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13656 n_53580_87640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13657 n_57000_87640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13658 n_65360_65240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13659 n_63460_62440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13660 n_63460_59640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13661 n_63460_56840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13662 n_68780_59640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13663 n_66880_59640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13664 n_70300_59640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13665 n_70300_56840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13666 n_71820_59640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13667 n_70300_65240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13668 n_68400_65240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13669 n_71820_68040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13670 n_73720_65240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13671 n_70300_70840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13672 n_67260_76440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13673 n_68780_76440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13674 n_65740_79240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13675 n_64600_79240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13676 n_57380_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13677 n_55100_79240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13678 n_58520_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13679 n_59660_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13680 n_56240_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13681 n_87400_62440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13682 n_88920_62440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13683 n_87020_59640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13684 n_85880_62440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13685 n_83220_65240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13686 n_83220_62440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13687 n_83220_68040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13688 n_84740_68040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13689 n_83600_70840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13690 n_83220_73640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13691 n_85880_73640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13692 n_83600_76440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13693 n_85500_76440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13694 n_85500_79240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13695 n_83600_79240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13696 n_85500_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13697 n_68780_82040 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13698 n_43320_65240 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13699 n_40280_62440 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13700 n_44460_56840 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13701 n_60040_59640 0 PWL(120000ps 0uA 120030ps 0uA 120031ps 30uA 120059ps 30uA 120060ps 0uA)
I13702 n_93480_79240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13703 n_91960_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13704 n_87020_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13705 n_93100_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13706 n_90440_62440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13707 n_83600_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13708 n_84740_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13709 n_56240_48440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13710 n_65740_45640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13711 n_61940_48440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13712 n_40280_54040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13713 n_40660_56840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13714 n_63840_45640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13715 n_93480_48440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13716 n_93480_54040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13717 n_92340_48440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13718 n_50920_48440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13719 n_63840_40040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13720 n_70300_40040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13721 n_91580_40040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13722 n_87020_40040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13723 n_42940_42840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13724 n_67260_40040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13725 n_60040_45640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13726 n_72200_40040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13727 n_79040_40040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13728 n_82080_48440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13729 n_77140_40040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13730 n_42180_73640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13731 n_40660_65240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13732 n_47500_40040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13733 n_89300_48440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13734 n_41800_68040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13735 n_52060_73640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13736 n_74860_40040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13737 n_80180_45640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13738 n_76760_42840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13739 n_71820_42840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13740 n_56620_45640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13741 n_66880_45640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13742 n_44840_45640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13743 n_87020_45640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13744 n_92720_40040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13745 n_68400_40040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13746 n_63460_42840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13747 n_51680_48440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13748 n_85120_48440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13749 n_92340_51240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13750 n_90440_48440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13751 n_64980_48440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13752 n_41420_54040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13753 n_47880_54040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13754 n_60040_48440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13755 n_64600_51240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13756 n_55100_54040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13757 n_81700_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13758 n_80180_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13759 n_90820_59640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13760 n_90060_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13761 n_85120_84840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13762 n_87400_84840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13763 n_91580_79240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13764 n_73340_51240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13765 n_71820_48440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13766 n_73340_48440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13767 n_68780_79240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13768 n_73720_54040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13769 n_87780_54040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13770 n_88920_51240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13771 n_83220_54040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13772 n_91200_54040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13773 n_92340_56840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13774 n_90820_65240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13775 n_88920_70840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13776 n_87400_65240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13777 n_87400_70840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13778 n_87400_76440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13779 n_92340_76440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13780 n_87780_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13781 n_82080_84840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13782 n_85880_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13783 n_83600_51240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13784 n_80560_51240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13785 n_84740_54040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13786 n_92720_59640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13787 n_77900_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13788 n_79040_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13789 n_79040_54040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13790 n_80560_54040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13791 n_82080_54040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13792 n_76760_56840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13793 n_79040_68040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13794 n_67260_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13795 n_65740_84840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13796 n_62320_82040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13797 n_65360_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13798 n_68780_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13799 n_71820_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13800 n_72200_84840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13801 n_85500_56840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13802 n_82080_59640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13803 n_85500_59640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13804 n_84740_65240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13805 n_83600_59640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13806 n_82080_65240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13807 n_82080_68040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13808 n_82080_70840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13809 n_80560_68040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13810 n_77140_70840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13811 n_81700_73640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13812 n_80560_73640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13813 n_78660_73640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13814 n_79040_70840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13815 n_80560_79240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13816 n_74860_84840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13817 n_74860_82040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13818 n_76760_82040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13819 n_60800_51240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13820 n_67260_51240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13821 n_71820_51240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13822 n_71820_54040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13823 n_53200_51240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13824 n_70300_51240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13825 n_68020_54040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13826 n_68780_51240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13827 n_59280_51240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13828 n_49780_54040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13829 n_41800_56840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13830 n_75240_54040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13831 n_66120_51240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13832 n_76380_51240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13833 n_79040_51240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13834 n_76760_48440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13835 n_87400_51240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13836 n_90820_51240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13837 n_85500_45640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13838 n_49400_48440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13839 n_50160_45640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13840 n_48260_48440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13841 n_61560_42840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13842 n_70300_42840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13843 n_89300_40040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13844 n_90440_45640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13845 n_85500_40040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13846 n_81700_40040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13847 n_46740_45640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13848 n_68780_45640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13849 n_82080_42840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13850 n_73720_42840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13851 n_58520_45640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13852 n_73720_45640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13853 n_76760_45640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13854 n_80560_48440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13855 n_73340_40040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13856 n_48640_59640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13857 n_49780_56840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13858 n_48260_62440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13859 n_48260_65240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13860 n_49780_62440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13861 n_59660_62440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13862 n_44840_73640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13863 n_50920_68040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13864 n_40280_59640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13865 n_56620_65240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13866 n_58520_65240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13867 n_60420_65240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13868 n_73720_62440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13869 n_63460_68040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13870 n_60040_73640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13871 n_76380_62440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13872 n_63080_82040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13873 n_75240_59640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13874 n_72200_62440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13875 n_61940_68040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13876 n_59660_70840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13877 n_53580_73640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13878 n_50920_73640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13879 n_48260_73640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13880 n_49780_76440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13881 n_50920_79240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13882 n_46360_79240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13883 n_58520_68040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13884 n_58520_73640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13885 n_70300_73640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13886 n_74100_68040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13887 n_75240_68040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13888 n_72960_68040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13889 n_68020_62440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13890 n_55480_48440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13891 n_40280_73640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13892 n_48260_76440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13893 n_47500_79240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13894 n_45600_84840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13895 n_48640_79240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13896 n_58520_70840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13897 n_49400_79240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13898 n_60040_76440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13899 n_60420_70840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13900 n_76760_73640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13901 n_60040_79240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13902 n_63080_79240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13903 n_70300_48440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13904 n_63080_76440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13905 n_49400_82040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13906 n_54720_84840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13907 n_65740_73640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13908 n_70300_76440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13909 n_47500_56840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13910 n_52820_79240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13911 n_41420_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13912 n_46740_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13913 n_43320_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13914 n_61940_84840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13915 n_52440_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13916 n_58140_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13917 n_55100_82040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13918 n_61940_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13919 n_42940_54040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13920 n_46740_51240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13921 n_41800_65240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13922 n_65360_59640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13923 n_66880_62440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13924 n_65360_54040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13925 n_63080_54040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13926 n_45220_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13927 n_59280_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13928 n_51680_84840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13929 n_60800_84840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13930 n_61180_82040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13931 n_54340_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13932 n_67260_82040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13933 n_65740_82040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13934 n_53580_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13935 n_58520_84840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13936 n_64600_84840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13937 n_57000_87640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13938 n_67260_65240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13939 n_63460_62440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13940 n_66880_59640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13941 n_70300_59640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13942 n_70300_62440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13943 n_71820_59640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13944 n_70300_65240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13945 n_68400_65240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13946 n_71820_68040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13947 n_70300_70840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13948 n_67260_76440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13949 n_68780_76440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13950 n_65740_79240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13951 n_53960_79240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13952 n_55100_79240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13953 n_56240_82040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13954 n_87400_62440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13955 n_88920_62440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13956 n_85880_62440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13957 n_83220_65240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13958 n_83220_62440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13959 n_83220_68040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13960 n_83600_70840 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13961 n_83220_73640 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13962 n_85500_82040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13963 n_68780_82040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13964 n_71060_82040 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13965 n_43320_65240 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13966 n_40280_62440 0 PWL(122000ps 0uA 122030ps 0uA 122031ps 30uA 122059ps 30uA 122060ps 0uA)
I13967 n_92340_54040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13968 n_90820_68040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13969 n_93480_79240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13970 n_93480_56840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13971 n_90440_62440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13972 n_93480_68040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13973 n_93480_73640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13974 n_93100_84840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13975 n_56240_48440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13976 n_61940_48440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13977 n_40280_54040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13978 n_44080_54040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13979 n_63840_45640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13980 n_79040_42840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13981 n_93480_48440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13982 n_93480_54040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13983 n_41800_42840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13984 n_50920_48440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13985 n_91580_40040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13986 n_87020_40040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13987 n_88160_40040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13988 n_40660_42840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13989 n_42940_42840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13990 n_40280_40040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13991 n_40280_48440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13992 n_60040_45640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13993 n_82080_48440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13994 n_43320_59640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13995 n_40660_65240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13996 n_41800_68040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13997 n_46740_59640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13998 n_80180_45640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I13999 n_56620_45640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14000 n_41420_48440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14001 n_41420_40040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14002 n_44840_45640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14003 n_43700_42840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14004 n_83600_40040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14005 n_87020_45640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14006 n_92720_40040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14007 n_51680_48440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14008 n_48260_45640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14009 n_92340_51240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14010 n_90440_48440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14011 n_78280_48440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14012 n_64980_48440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14013 n_49020_51240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14014 n_47880_54040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14015 n_60040_48440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14016 n_55100_54040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14017 n_90820_84840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14018 n_90440_73640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14019 n_92340_65240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14020 n_90820_59640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14021 n_88920_56840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14022 n_91580_79240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14023 n_88540_68040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14024 n_89300_54040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14025 n_87780_54040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14026 n_83220_54040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14027 n_91200_54040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14028 n_92340_56840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14029 n_90820_65240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14030 n_88920_70840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14031 n_87400_70840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14032 n_87400_76440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14033 n_92340_76440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14034 n_87780_87640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14035 n_88920_82040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14036 n_83600_51240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14037 n_80560_51240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14038 n_84740_54040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14039 n_90820_56840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14040 n_92720_59640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14041 n_91960_68040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14042 n_92340_73640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14043 n_90820_82040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14044 n_82080_54040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14045 n_80560_56840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14046 n_80180_59640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14047 n_78660_56840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14048 n_83600_56840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14049 n_76380_54040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14050 n_76760_65240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14051 n_76760_56840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14052 n_76380_68040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14053 n_78660_65240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14054 n_77900_68040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14055 n_76000_70840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14056 n_79040_68040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14057 n_78280_70840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14058 n_75240_73640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14059 n_73720_70840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14060 n_73720_79240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14061 n_70300_79240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14062 n_67260_84840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14063 n_65740_84840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14064 n_62320_82040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14065 n_68780_84840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14066 n_71820_87640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14067 n_70300_87640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14068 n_85500_56840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14069 n_87400_48440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14070 n_82080_59640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14071 n_85500_59640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14072 n_84740_65240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14073 n_83600_59640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14074 n_82080_65240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14075 n_82080_68040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14076 n_87400_68040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14077 n_82080_70840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14078 n_77140_70840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14079 n_81700_73640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14080 n_80560_70840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14081 n_80560_73640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14082 n_78660_73640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14083 n_79040_70840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14084 n_78280_82040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14085 n_76760_79240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14086 n_76760_84840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14087 n_76380_87640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14088 n_60800_51240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14089 n_67260_51240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14090 n_71820_51240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14091 n_71820_54040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14092 n_53200_51240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14093 n_70300_51240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14094 n_68020_54040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14095 n_56620_51240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14096 n_68780_51240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14097 n_59280_51240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14098 n_49780_54040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14099 n_47880_51240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14100 n_70300_54040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14101 n_61560_54040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14102 n_66120_51240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14103 n_79040_51240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14104 n_87400_51240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14105 n_90820_51240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14106 n_49400_48440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14107 n_53200_48440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14108 n_92720_42840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14109 n_90440_45640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14110 n_85500_40040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14111 n_45220_42840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14112 n_46740_45640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14113 n_43320_40040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14114 n_42940_48440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14115 n_53200_45640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14116 n_82080_45640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14117 n_58900_48440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14118 n_49780_56840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14119 n_48260_62440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14120 n_48260_65240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14121 n_49780_62440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14122 n_59660_62440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14123 n_44840_73640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14124 n_50920_68040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14125 n_56620_65240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14126 n_61560_62440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14127 n_61560_65240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14128 n_59660_68040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14129 n_60800_68040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14130 n_60040_73640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14131 n_63080_65240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14132 n_75240_59640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14133 n_73340_59640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14134 n_61940_68040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14135 n_59660_70840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14136 n_49400_73640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14137 n_55860_68040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14138 n_46740_73640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14139 n_46360_76440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14140 n_40660_76440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14141 n_48260_73640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14142 n_40660_70840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14143 n_49780_76440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14144 n_50920_79240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14145 n_58520_73640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14146 n_70300_73640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14147 n_66880_73640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14148 n_58140_79240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14149 n_63460_70840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14150 n_74100_68040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14151 n_65360_70840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14152 n_68780_68040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14153 n_75240_68040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14154 n_72960_68040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14155 n_48260_76440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14156 n_47500_79240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14157 n_48640_79240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14158 n_58520_70840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14159 n_60040_76440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14160 n_60420_70840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14161 n_76760_73640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14162 n_56620_79240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14163 n_52060_82040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14164 n_68400_73640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14165 n_40660_79240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14166 n_40280_82040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14167 n_43700_79240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14168 n_40280_87640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14169 n_57380_76440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14170 n_50920_82040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14171 n_53580_82040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14172 n_47500_56840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14173 n_40280_84840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14174 n_41420_87640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14175 n_46740_87640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14176 n_46740_84840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14177 n_49400_84840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14178 n_61940_87640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14179 n_43320_68040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14180 n_43320_76440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14181 n_44080_82040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14182 n_65360_62440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14183 n_66880_62440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14184 n_65360_56840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14185 n_68780_56840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14186 n_54340_76440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14187 n_56240_76440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14188 n_65360_65240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14189 n_67260_65240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14190 n_60040_54040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14191 n_67260_56840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14192 n_70300_59640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14193 n_70300_62440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14194 n_71820_59640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14195 n_70300_65240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14196 n_68400_65240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14197 n_73720_65240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14198 n_64600_79240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14199 n_53960_79240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14200 n_57380_82040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14201 n_58520_82040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14202 n_59660_82040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14203 n_87400_62440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14204 n_88920_62440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14205 n_88160_59640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14206 n_85880_62440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14207 n_83220_65240 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14208 n_83220_62440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14209 n_83220_68040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14210 n_83600_70840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14211 n_85500_70840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14212 n_84740_73640 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14213 n_83600_76440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14214 n_85500_76440 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14215 n_87400_82040 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14216 n_44460_56840 0 PWL(124000ps 0uA 124030ps 0uA 124031ps 30uA 124059ps 30uA 124060ps 0uA)
I14217 n_91200_70840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14218 n_93100_87640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14219 n_93480_68040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14220 n_93480_73640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14221 n_93480_76440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14222 n_84740_87640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14223 n_65740_45640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14224 n_61940_48440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14225 n_40280_54040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14226 n_44080_54040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14227 n_40660_56840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14228 n_63840_45640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14229 n_79040_42840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14230 n_41800_42840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14231 n_63840_40040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14232 n_91580_40040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14233 n_87020_40040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14234 n_40660_42840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14235 n_56620_40040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14236 n_67260_40040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14237 n_93480_45640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14238 n_80560_40040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14239 n_46360_40040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14240 n_72200_40040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14241 n_82080_48440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14242 n_77140_40040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14243 n_40660_45640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14244 n_40660_51240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14245 n_50160_59640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14246 n_42180_73640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14247 n_45600_68040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14248 n_43320_62440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14249 n_40660_65240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14250 n_41800_68040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14251 n_44460_62440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14252 n_47500_68040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14253 n_52060_73640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14254 n_51300_59640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14255 n_44840_51240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14256 n_45220_48440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14257 n_74860_40040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14258 n_80180_45640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14259 n_71820_42840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14260 n_49400_40040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14261 n_80180_42840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14262 n_88920_45640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14263 n_66880_45640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14264 n_57760_40040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14265 n_43700_42840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14266 n_87020_45640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14267 n_92720_40040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14268 n_63460_42840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14269 n_48260_45640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14270 n_78280_48440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14271 n_64980_48440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14272 n_41420_54040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14273 n_49020_51240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14274 n_47880_54040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14275 n_60040_48440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14276 n_64600_51240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14277 n_81700_87640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14278 n_90440_76440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14279 n_90440_73640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14280 n_92340_65240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14281 n_90060_87640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14282 n_87400_73640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14283 n_87400_76440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14284 n_85880_87640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14285 n_91960_68040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14286 n_92340_73640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14287 n_90060_79240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14288 n_79040_87640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14289 n_78660_56840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14290 n_83600_56840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14291 n_76380_54040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14292 n_80940_62440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14293 n_76760_56840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14294 n_76380_68040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14295 n_78280_70840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14296 n_75240_76440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14297 n_73720_73640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14298 n_88920_79240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14299 n_62320_82040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14300 n_68780_87640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14301 n_68780_84840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14302 n_86260_54040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14303 n_85500_59640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14304 n_80560_70840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14305 n_80560_73640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14306 n_78280_82040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14307 n_76760_79240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14308 n_76760_84840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14309 n_76380_87640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14310 n_74860_84840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14311 n_60800_51240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14312 n_67260_51240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14313 n_71820_51240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14314 n_71820_54040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14315 n_53200_51240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14316 n_70300_51240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14317 n_56620_51240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14318 n_59280_51240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14319 n_49780_54040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14320 n_47880_51240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14321 n_52060_51240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14322 n_70300_54040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14323 n_61560_54040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14324 n_66120_51240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14325 n_79040_51240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14326 n_49400_48440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14327 n_65360_42840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14328 n_92720_42840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14329 n_90440_45640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14330 n_45220_42840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14331 n_61560_40040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14332 n_68020_48440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14333 n_88920_42840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14334 n_82080_42840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14335 n_51300_40040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14336 n_73720_45640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14337 n_82080_45640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14338 n_73340_40040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14339 n_44080_48440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14340 n_43320_51240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14341 n_57000_54040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14342 n_52060_54040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14343 n_48260_65240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14344 n_59660_62440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14345 n_50920_68040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14346 n_72200_56840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14347 n_53580_59640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14348 n_53580_62440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14349 n_52060_65240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14350 n_49400_65240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14351 n_56620_65240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14352 n_61560_62440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14353 n_61560_65240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14354 n_59660_68040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14355 n_60800_68040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14356 n_63460_68040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14357 n_63080_65240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14358 n_76380_59640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14359 n_55100_56840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14360 n_55100_70840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14361 n_53580_70840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14362 n_50920_70840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14363 n_50920_73640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14364 n_49400_73640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14365 n_55860_68040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14366 n_49780_76440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14367 n_50920_79240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14368 n_58520_68040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14369 n_70300_73640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14370 n_56620_73640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14371 n_66880_73640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14372 n_63460_70840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14373 n_65360_70840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14374 n_68780_68040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14375 n_72960_68040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14376 n_68780_70840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14377 n_47500_79240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14378 n_48640_79240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14379 n_60040_76440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14380 n_63080_73640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14381 n_76760_73640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14382 n_61560_79240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14383 n_65740_76440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14384 n_68400_73640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14385 n_58140_51240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14386 n_46360_68040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14387 n_44840_70840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14388 n_43320_70840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14389 n_41800_70840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14390 n_40660_79240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14391 n_43700_79240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14392 n_57380_76440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14393 n_70300_76440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14394 n_52820_79240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14395 n_44080_59640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14396 n_42940_82040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14397 n_42940_84840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14398 n_42940_54040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14399 n_46740_51240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14400 n_43320_68040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14401 n_43320_76440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14402 n_44080_82040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14403 n_65360_62440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14404 n_66880_62440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14405 n_65360_65240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14406 n_67260_65240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14407 n_63460_59640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14408 n_63460_56840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14409 n_60040_54040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14410 n_70300_59640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14411 n_70300_56840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14412 n_71820_59640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14413 n_71820_65240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14414 n_71820_68040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14415 n_70300_70840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14416 n_71820_70840 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14417 n_67260_76440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14418 n_65740_79240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14419 n_64600_79240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14420 n_57380_82040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14421 n_58520_82040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14422 n_56240_82040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14423 n_87400_62440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14424 n_87020_59640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14425 n_88160_59640 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14426 n_85880_62440 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14427 n_83220_65240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14428 n_83220_68040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14429 n_84740_68040 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14430 n_85500_79240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14431 n_83600_79240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14432 n_43320_65240 0 PWL(126000ps 0uA 126030ps 0uA 126031ps 30uA 126059ps 30uA 126060ps 0uA)
I14433 n_90820_68040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14434 n_91200_70840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14435 n_93480_79240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14436 n_93480_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14437 n_93100_84840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14438 n_54720_48440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14439 n_61940_48440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14440 n_40660_56840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14441 n_79040_42840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14442 n_92340_48440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14443 n_50920_48440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14444 n_91580_40040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14445 n_40660_42840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14446 n_67260_40040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14447 n_90440_40040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14448 n_93480_45640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14449 n_46360_40040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14450 n_60040_45640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14451 n_72200_40040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14452 n_82080_48440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14453 n_55100_40040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14454 n_43320_59640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14455 n_50160_59640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14456 n_42180_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14457 n_45600_68040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14458 n_43320_62440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14459 n_44460_62440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14460 n_47500_68040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14461 n_52060_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14462 n_51300_59640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14463 n_46740_59640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14464 n_54720_42840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14465 n_80180_45640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14466 n_71820_42840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14467 n_56620_45640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14468 n_49400_40040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14469 n_88920_45640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14470 n_83600_42840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14471 n_66880_45640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14472 n_43700_42840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14473 n_92720_40040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14474 n_51680_48440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14475 n_85120_48440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14476 n_78280_48440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14477 n_41420_54040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14478 n_60040_48440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14479 n_54720_51240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14480 n_90820_84840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14481 n_90440_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14482 n_91580_79240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14483 n_87400_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14484 n_88540_68040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14485 n_87400_65240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14486 n_87400_76440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14487 n_92340_76440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14488 n_92340_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14489 n_90820_82040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14490 n_76760_65240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14491 n_80940_62440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14492 n_76760_56840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14493 n_78660_65240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14494 n_77900_68040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14495 n_76000_70840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14496 n_75240_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14497 n_75240_76440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14498 n_73720_79240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14499 n_73720_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14500 n_70300_79240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14501 n_67260_84840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14502 n_65740_84840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14503 n_70300_87640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14504 n_85500_59640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14505 n_87400_68040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14506 n_80560_68040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14507 n_81700_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14508 n_80560_70840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14509 n_80560_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14510 n_81700_76440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14511 n_76760_76440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14512 n_72200_76440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14513 n_70300_51240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14514 n_61940_51240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14515 n_52060_51240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14516 n_79040_51240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14517 n_83600_48440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14518 n_53200_48440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14519 n_92720_42840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14520 n_45220_42840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14521 n_68020_48440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14522 n_85500_42840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14523 n_88920_42840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14524 n_51300_40040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14525 n_53200_45640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14526 n_73720_45640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14527 n_82080_45640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14528 n_53200_42840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14529 n_58900_48440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14530 n_57000_54040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14531 n_49780_56840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14532 n_48260_62440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14533 n_49780_62440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14534 n_44840_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14535 n_72200_56840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14536 n_53580_59640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14537 n_53580_62440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14538 n_52060_65240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14539 n_49400_65240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14540 n_63460_68040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14541 n_60040_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14542 n_76380_59640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14543 n_61940_68040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14544 n_59660_70840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14545 n_55100_56840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14546 n_55100_70840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14547 n_53580_70840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14548 n_50920_70840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14549 n_50920_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14550 n_46740_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14551 n_46360_76440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14552 n_40660_76440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14553 n_48260_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14554 n_40660_70840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14555 n_58520_68040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14556 n_61560_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14557 n_70300_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14558 n_56620_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14559 n_66880_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14560 n_58140_79240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14561 n_74100_68040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14562 n_75240_68040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14563 n_55480_48440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14564 n_68780_70840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14565 n_48260_76440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14566 n_58520_70840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14567 n_60420_70840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14568 n_76760_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14569 n_60040_79240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14570 n_63080_79240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14571 n_61560_79240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14572 n_52060_82040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14573 n_68400_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14574 n_58140_51240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14575 n_46360_68040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14576 n_44840_70840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14577 n_43320_70840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14578 n_41800_70840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14579 n_40280_82040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14580 n_40280_87640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14581 n_57380_76440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14582 n_67260_79240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14583 n_80560_76440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14584 n_50920_82040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14585 n_53580_82040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14586 n_47500_56840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14587 n_52820_79240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14588 n_44080_59640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14589 n_42940_82040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14590 n_42940_84840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14591 n_40280_84840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14592 n_41420_87640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14593 n_46740_87640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14594 n_46740_84840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14595 n_49400_84840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14596 n_61940_87640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14597 n_42940_54040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14598 n_65360_56840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14599 n_68780_56840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14600 n_54340_76440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14601 n_56240_76440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14602 n_63460_59640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14603 n_63460_56840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14604 n_60040_54040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14605 n_67260_56840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14606 n_66880_59640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14607 n_70300_59640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14608 n_70300_56840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14609 n_71820_59640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14610 n_71820_65240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14611 n_71820_68040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14612 n_70300_70840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14613 n_71820_70840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14614 n_67260_76440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14615 n_65740_79240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14616 n_64600_79240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14617 n_53960_79240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14618 n_64600_76440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14619 n_59660_82040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14620 n_84740_68040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14621 n_83600_70840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14622 n_85500_70840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14623 n_84740_73640 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14624 n_83600_76440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14625 n_85500_76440 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14626 n_85500_79240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14627 n_87400_82040 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14628 n_83600_79240 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14629 n_44460_56840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14630 n_60040_56840 0 PWL(128000ps 0uA 128030ps 0uA 128031ps 30uA 128059ps 30uA 128060ps 0uA)
I14631 n_91200_70840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14632 n_93100_87640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14633 n_93480_73640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14634 n_93480_76440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14635 n_93100_84840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14636 n_84740_87640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14637 n_65740_40040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14638 n_40280_54040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14639 n_40660_56840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14640 n_63840_45640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14641 n_79040_42840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14642 n_92340_48440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14643 n_48640_40040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14644 n_50920_48440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14645 n_88160_40040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14646 n_52440_40040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14647 n_42940_42840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14648 n_56620_40040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14649 n_93480_45640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14650 n_40280_48440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14651 n_79040_40040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14652 n_82080_48440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14653 n_55100_40040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14654 n_40660_45640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14655 n_43320_59640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14656 n_50160_59640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14657 n_42180_73640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14658 n_44460_68040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14659 n_45600_68040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14660 n_43320_62440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14661 n_44460_62440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14662 n_47500_68040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14663 n_46740_65240 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14664 n_52060_73640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14665 n_51300_59640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14666 n_46740_59640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14667 n_45220_48440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14668 n_54720_42840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14669 n_80180_45640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14670 n_76760_42840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14671 n_41420_48440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14672 n_88920_45640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14673 n_57760_40040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14674 n_44840_45640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14675 n_51680_42840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14676 n_83600_40040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14677 n_51680_48440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14678 n_47880_42840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14679 n_85120_48440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14680 n_78280_48440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14681 n_64980_48440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14682 n_41420_54040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14683 n_47880_54040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14684 n_63080_51240 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14685 n_81700_87640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14686 n_90820_84840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14687 n_90440_76440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14688 n_90440_73640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14689 n_90060_87640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14690 n_87400_73640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14691 n_87400_76440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14692 n_85880_87640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14693 n_92340_73640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14694 n_90060_79240 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14695 n_90820_82040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14696 n_79040_87640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14697 n_83600_56840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14698 n_76380_54040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14699 n_76760_65240 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14700 n_80940_62440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14701 n_76760_56840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14702 n_78660_65240 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14703 n_77900_68040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14704 n_76000_70840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14705 n_75240_73640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14706 n_73720_79240 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14707 n_73720_73640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14708 n_88920_79240 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14709 n_67260_87640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14710 n_65740_84840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14711 n_65360_87640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14712 n_70300_87640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14713 n_73720_82040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14714 n_86260_54040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14715 n_85500_59640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14716 n_82080_70840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14717 n_80560_70840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14718 n_80560_73640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14719 n_81700_76440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14720 n_78660_73640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14721 n_78660_76440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14722 n_78660_79240 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14723 n_72200_76440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14724 n_78280_82040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14725 n_80180_82040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14726 n_76760_84840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14727 n_76380_87640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14728 n_74860_84840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14729 n_67260_51240 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14730 n_71820_51240 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14731 n_71820_54040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14732 n_59280_51240 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14733 n_61940_51240 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14734 n_49780_54040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14735 n_41800_56840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14736 n_70300_54040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14737 n_61560_54040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14738 n_66120_51240 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14739 n_79040_51240 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14740 n_83600_48440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14741 n_51680_45640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14742 n_53200_48440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14743 n_85500_40040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14744 n_50540_42840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14745 n_46740_45640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14746 n_61560_40040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14747 n_88920_42840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14748 n_42940_48440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14749 n_76760_45640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14750 n_82080_45640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14751 n_53200_42840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14752 n_44080_48440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14753 n_58900_48440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14754 n_57000_54040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14755 n_49780_56840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14756 n_48260_62440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14757 n_49780_62440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14758 n_44840_73640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14759 n_53580_59640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14760 n_53580_62440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14761 n_52060_65240 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14762 n_49400_65240 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14763 n_76380_59640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14764 n_69160_62440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14765 n_55100_70840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14766 n_53580_70840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14767 n_50920_70840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14768 n_50920_73640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14769 n_46740_73640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14770 n_40660_76440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14771 n_40660_70840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14772 n_61560_73640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14773 n_58520_73640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14774 n_70300_73640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14775 n_66880_73640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14776 n_53580_65240 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14777 n_53580_68040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14778 n_49400_70840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14779 n_46740_70840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14780 n_63080_73640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14781 n_76760_73640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14782 n_52060_82040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14783 n_65740_76440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14784 n_68400_73640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14785 n_70300_48440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14786 n_46360_68040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14787 n_44840_70840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14788 n_43320_70840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14789 n_41800_70840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14790 n_40280_82040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14791 n_40280_87640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14792 n_50920_82040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14793 n_53580_82040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14794 n_70300_76440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14795 n_47500_56840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14796 n_44080_59640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14797 n_42940_82040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14798 n_42940_84840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14799 n_40280_84840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14800 n_41420_87640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14801 n_46740_87640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14802 n_46740_84840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14803 n_49400_84840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14804 n_61940_87640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14805 n_42940_54040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14806 n_46740_51240 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14807 n_65360_56840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14808 n_68780_56840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14809 n_54340_76440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14810 n_56240_76440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14811 n_67260_56840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14812 n_66880_59640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14813 n_71820_59640 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14814 n_68400_65240 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14815 n_71820_65240 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14816 n_71820_68040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14817 n_70300_70840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14818 n_67260_76440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14819 n_68780_76440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14820 n_57380_82040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14821 n_64600_76440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14822 n_58520_82040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14823 n_59660_82040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14824 n_56240_82040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14825 n_56620_84840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14826 n_81700_79240 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14827 n_85500_76440 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14828 n_87400_82040 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14829 n_44460_56840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
I14830 n_60040_56840 0 PWL(130000ps 0uA 130030ps 0uA 130031ps 30uA 130059ps 30uA 130060ps 0uA)
.tran 1ps 134000ps
.control
run
* calculate minimum value of voltage at each node:
let min_40280_40040 = minimum(v(n_40280_40040))
let min_40280_42840 = minimum(v(n_40280_42840))
let min_40280_45640 = minimum(v(n_40280_45640))
let min_40280_48440 = minimum(v(n_40280_48440))
let min_40280_51240 = minimum(v(n_40280_51240))
let min_40280_54040 = minimum(v(n_40280_54040))
let min_40280_56840 = minimum(v(n_40280_56840))
let min_40280_59640 = minimum(v(n_40280_59640))
let min_40280_62440 = minimum(v(n_40280_62440))
let min_40280_65240 = minimum(v(n_40280_65240))
let min_40280_68040 = minimum(v(n_40280_68040))
let min_40280_70840 = minimum(v(n_40280_70840))
let min_40280_73640 = minimum(v(n_40280_73640))
let min_40280_76440 = minimum(v(n_40280_76440))
let min_40280_79240 = minimum(v(n_40280_79240))
let min_40280_82040 = minimum(v(n_40280_82040))
let min_40280_84840 = minimum(v(n_40280_84840))
let min_40280_87640 = minimum(v(n_40280_87640))
let min_40660_40040 = minimum(v(n_40660_40040))
let min_40660_42840 = minimum(v(n_40660_42840))
let min_40660_45640 = minimum(v(n_40660_45640))
let min_40660_48440 = minimum(v(n_40660_48440))
let min_40660_51240 = minimum(v(n_40660_51240))
let min_40660_54040 = minimum(v(n_40660_54040))
let min_40660_56840 = minimum(v(n_40660_56840))
let min_40660_59640 = minimum(v(n_40660_59640))
let min_40660_62440 = minimum(v(n_40660_62440))
let min_40660_65240 = minimum(v(n_40660_65240))
let min_40660_68040 = minimum(v(n_40660_68040))
let min_40660_70840 = minimum(v(n_40660_70840))
let min_40660_73640 = minimum(v(n_40660_73640))
let min_40660_76440 = minimum(v(n_40660_76440))
let min_40660_79240 = minimum(v(n_40660_79240))
let min_40660_82040 = minimum(v(n_40660_82040))
let min_40660_84840 = minimum(v(n_40660_84840))
let min_40660_87640 = minimum(v(n_40660_87640))
let min_41420_40040 = minimum(v(n_41420_40040))
let min_41420_42840 = minimum(v(n_41420_42840))
let min_41420_45640 = minimum(v(n_41420_45640))
let min_41420_48440 = minimum(v(n_41420_48440))
let min_41420_51240 = minimum(v(n_41420_51240))
let min_41420_54040 = minimum(v(n_41420_54040))
let min_41420_56840 = minimum(v(n_41420_56840))
let min_41420_59640 = minimum(v(n_41420_59640))
let min_41420_62440 = minimum(v(n_41420_62440))
let min_41420_65240 = minimum(v(n_41420_65240))
let min_41420_68040 = minimum(v(n_41420_68040))
let min_41420_70840 = minimum(v(n_41420_70840))
let min_41420_73640 = minimum(v(n_41420_73640))
let min_41420_76440 = minimum(v(n_41420_76440))
let min_41420_79240 = minimum(v(n_41420_79240))
let min_41420_82040 = minimum(v(n_41420_82040))
let min_41420_84840 = minimum(v(n_41420_84840))
let min_41420_87640 = minimum(v(n_41420_87640))
let min_41800_40040 = minimum(v(n_41800_40040))
let min_41800_42840 = minimum(v(n_41800_42840))
let min_41800_45640 = minimum(v(n_41800_45640))
let min_41800_48440 = minimum(v(n_41800_48440))
let min_41800_51240 = minimum(v(n_41800_51240))
let min_41800_54040 = minimum(v(n_41800_54040))
let min_41800_56840 = minimum(v(n_41800_56840))
let min_41800_59640 = minimum(v(n_41800_59640))
let min_41800_62440 = minimum(v(n_41800_62440))
let min_41800_65240 = minimum(v(n_41800_65240))
let min_41800_68040 = minimum(v(n_41800_68040))
let min_41800_70840 = minimum(v(n_41800_70840))
let min_41800_73640 = minimum(v(n_41800_73640))
let min_41800_76440 = minimum(v(n_41800_76440))
let min_41800_79240 = minimum(v(n_41800_79240))
let min_41800_82040 = minimum(v(n_41800_82040))
let min_41800_84840 = minimum(v(n_41800_84840))
let min_41800_87640 = minimum(v(n_41800_87640))
let min_42180_40040 = minimum(v(n_42180_40040))
let min_42180_42840 = minimum(v(n_42180_42840))
let min_42180_45640 = minimum(v(n_42180_45640))
let min_42180_48440 = minimum(v(n_42180_48440))
let min_42180_51240 = minimum(v(n_42180_51240))
let min_42180_54040 = minimum(v(n_42180_54040))
let min_42180_56840 = minimum(v(n_42180_56840))
let min_42180_59640 = minimum(v(n_42180_59640))
let min_42180_62440 = minimum(v(n_42180_62440))
let min_42180_65240 = minimum(v(n_42180_65240))
let min_42180_68040 = minimum(v(n_42180_68040))
let min_42180_70840 = minimum(v(n_42180_70840))
let min_42180_73640 = minimum(v(n_42180_73640))
let min_42180_76440 = minimum(v(n_42180_76440))
let min_42180_79240 = minimum(v(n_42180_79240))
let min_42180_82040 = minimum(v(n_42180_82040))
let min_42180_84840 = minimum(v(n_42180_84840))
let min_42180_87640 = minimum(v(n_42180_87640))
let min_42940_40040 = minimum(v(n_42940_40040))
let min_42940_42840 = minimum(v(n_42940_42840))
let min_42940_45640 = minimum(v(n_42940_45640))
let min_42940_48440 = minimum(v(n_42940_48440))
let min_42940_51240 = minimum(v(n_42940_51240))
let min_42940_54040 = minimum(v(n_42940_54040))
let min_42940_56840 = minimum(v(n_42940_56840))
let min_42940_59640 = minimum(v(n_42940_59640))
let min_42940_62440 = minimum(v(n_42940_62440))
let min_42940_65240 = minimum(v(n_42940_65240))
let min_42940_68040 = minimum(v(n_42940_68040))
let min_42940_70840 = minimum(v(n_42940_70840))
let min_42940_73640 = minimum(v(n_42940_73640))
let min_42940_76440 = minimum(v(n_42940_76440))
let min_42940_79240 = minimum(v(n_42940_79240))
let min_42940_82040 = minimum(v(n_42940_82040))
let min_42940_84840 = minimum(v(n_42940_84840))
let min_42940_87640 = minimum(v(n_42940_87640))
let min_43320_40040 = minimum(v(n_43320_40040))
let min_43320_42840 = minimum(v(n_43320_42840))
let min_43320_45640 = minimum(v(n_43320_45640))
let min_43320_48440 = minimum(v(n_43320_48440))
let min_43320_51240 = minimum(v(n_43320_51240))
let min_43320_54040 = minimum(v(n_43320_54040))
let min_43320_56840 = minimum(v(n_43320_56840))
let min_43320_59640 = minimum(v(n_43320_59640))
let min_43320_62440 = minimum(v(n_43320_62440))
let min_43320_65240 = minimum(v(n_43320_65240))
let min_43320_68040 = minimum(v(n_43320_68040))
let min_43320_70840 = minimum(v(n_43320_70840))
let min_43320_73640 = minimum(v(n_43320_73640))
let min_43320_76440 = minimum(v(n_43320_76440))
let min_43320_79240 = minimum(v(n_43320_79240))
let min_43320_82040 = minimum(v(n_43320_82040))
let min_43320_84840 = minimum(v(n_43320_84840))
let min_43320_87640 = minimum(v(n_43320_87640))
let min_43700_40040 = minimum(v(n_43700_40040))
let min_43700_42840 = minimum(v(n_43700_42840))
let min_43700_45640 = minimum(v(n_43700_45640))
let min_43700_48440 = minimum(v(n_43700_48440))
let min_43700_51240 = minimum(v(n_43700_51240))
let min_43700_54040 = minimum(v(n_43700_54040))
let min_43700_56840 = minimum(v(n_43700_56840))
let min_43700_59640 = minimum(v(n_43700_59640))
let min_43700_62440 = minimum(v(n_43700_62440))
let min_43700_65240 = minimum(v(n_43700_65240))
let min_43700_68040 = minimum(v(n_43700_68040))
let min_43700_70840 = minimum(v(n_43700_70840))
let min_43700_73640 = minimum(v(n_43700_73640))
let min_43700_76440 = minimum(v(n_43700_76440))
let min_43700_79240 = minimum(v(n_43700_79240))
let min_43700_82040 = minimum(v(n_43700_82040))
let min_43700_84840 = minimum(v(n_43700_84840))
let min_43700_87640 = minimum(v(n_43700_87640))
let min_44080_40040 = minimum(v(n_44080_40040))
let min_44080_42840 = minimum(v(n_44080_42840))
let min_44080_45640 = minimum(v(n_44080_45640))
let min_44080_48440 = minimum(v(n_44080_48440))
let min_44080_51240 = minimum(v(n_44080_51240))
let min_44080_54040 = minimum(v(n_44080_54040))
let min_44080_56840 = minimum(v(n_44080_56840))
let min_44080_59640 = minimum(v(n_44080_59640))
let min_44080_62440 = minimum(v(n_44080_62440))
let min_44080_65240 = minimum(v(n_44080_65240))
let min_44080_68040 = minimum(v(n_44080_68040))
let min_44080_70840 = minimum(v(n_44080_70840))
let min_44080_73640 = minimum(v(n_44080_73640))
let min_44080_76440 = minimum(v(n_44080_76440))
let min_44080_79240 = minimum(v(n_44080_79240))
let min_44080_82040 = minimum(v(n_44080_82040))
let min_44080_84840 = minimum(v(n_44080_84840))
let min_44080_87640 = minimum(v(n_44080_87640))
let min_44460_40040 = minimum(v(n_44460_40040))
let min_44460_42840 = minimum(v(n_44460_42840))
let min_44460_45640 = minimum(v(n_44460_45640))
let min_44460_48440 = minimum(v(n_44460_48440))
let min_44460_51240 = minimum(v(n_44460_51240))
let min_44460_54040 = minimum(v(n_44460_54040))
let min_44460_56840 = minimum(v(n_44460_56840))
let min_44460_59640 = minimum(v(n_44460_59640))
let min_44460_62440 = minimum(v(n_44460_62440))
let min_44460_65240 = minimum(v(n_44460_65240))
let min_44460_68040 = minimum(v(n_44460_68040))
let min_44460_70840 = minimum(v(n_44460_70840))
let min_44460_73640 = minimum(v(n_44460_73640))
let min_44460_76440 = minimum(v(n_44460_76440))
let min_44460_79240 = minimum(v(n_44460_79240))
let min_44460_82040 = minimum(v(n_44460_82040))
let min_44460_84840 = minimum(v(n_44460_84840))
let min_44460_87640 = minimum(v(n_44460_87640))
let min_44840_40040 = minimum(v(n_44840_40040))
let min_44840_42840 = minimum(v(n_44840_42840))
let min_44840_45640 = minimum(v(n_44840_45640))
let min_44840_48440 = minimum(v(n_44840_48440))
let min_44840_51240 = minimum(v(n_44840_51240))
let min_44840_54040 = minimum(v(n_44840_54040))
let min_44840_56840 = minimum(v(n_44840_56840))
let min_44840_59640 = minimum(v(n_44840_59640))
let min_44840_62440 = minimum(v(n_44840_62440))
let min_44840_65240 = minimum(v(n_44840_65240))
let min_44840_68040 = minimum(v(n_44840_68040))
let min_44840_70840 = minimum(v(n_44840_70840))
let min_44840_73640 = minimum(v(n_44840_73640))
let min_44840_76440 = minimum(v(n_44840_76440))
let min_44840_79240 = minimum(v(n_44840_79240))
let min_44840_82040 = minimum(v(n_44840_82040))
let min_44840_84840 = minimum(v(n_44840_84840))
let min_44840_87640 = minimum(v(n_44840_87640))
let min_45220_40040 = minimum(v(n_45220_40040))
let min_45220_42840 = minimum(v(n_45220_42840))
let min_45220_45640 = minimum(v(n_45220_45640))
let min_45220_48440 = minimum(v(n_45220_48440))
let min_45220_51240 = minimum(v(n_45220_51240))
let min_45220_54040 = minimum(v(n_45220_54040))
let min_45220_56840 = minimum(v(n_45220_56840))
let min_45220_59640 = minimum(v(n_45220_59640))
let min_45220_62440 = minimum(v(n_45220_62440))
let min_45220_65240 = minimum(v(n_45220_65240))
let min_45220_68040 = minimum(v(n_45220_68040))
let min_45220_70840 = minimum(v(n_45220_70840))
let min_45220_73640 = minimum(v(n_45220_73640))
let min_45220_76440 = minimum(v(n_45220_76440))
let min_45220_79240 = minimum(v(n_45220_79240))
let min_45220_82040 = minimum(v(n_45220_82040))
let min_45220_84840 = minimum(v(n_45220_84840))
let min_45220_87640 = minimum(v(n_45220_87640))
let min_45600_40040 = minimum(v(n_45600_40040))
let min_45600_42840 = minimum(v(n_45600_42840))
let min_45600_45640 = minimum(v(n_45600_45640))
let min_45600_48440 = minimum(v(n_45600_48440))
let min_45600_51240 = minimum(v(n_45600_51240))
let min_45600_54040 = minimum(v(n_45600_54040))
let min_45600_56840 = minimum(v(n_45600_56840))
let min_45600_59640 = minimum(v(n_45600_59640))
let min_45600_62440 = minimum(v(n_45600_62440))
let min_45600_65240 = minimum(v(n_45600_65240))
let min_45600_68040 = minimum(v(n_45600_68040))
let min_45600_70840 = minimum(v(n_45600_70840))
let min_45600_73640 = minimum(v(n_45600_73640))
let min_45600_76440 = minimum(v(n_45600_76440))
let min_45600_79240 = minimum(v(n_45600_79240))
let min_45600_82040 = minimum(v(n_45600_82040))
let min_45600_84840 = minimum(v(n_45600_84840))
let min_45600_87640 = minimum(v(n_45600_87640))
let min_46360_40040 = minimum(v(n_46360_40040))
let min_46360_42840 = minimum(v(n_46360_42840))
let min_46360_45640 = minimum(v(n_46360_45640))
let min_46360_48440 = minimum(v(n_46360_48440))
let min_46360_51240 = minimum(v(n_46360_51240))
let min_46360_54040 = minimum(v(n_46360_54040))
let min_46360_56840 = minimum(v(n_46360_56840))
let min_46360_59640 = minimum(v(n_46360_59640))
let min_46360_62440 = minimum(v(n_46360_62440))
let min_46360_65240 = minimum(v(n_46360_65240))
let min_46360_68040 = minimum(v(n_46360_68040))
let min_46360_70840 = minimum(v(n_46360_70840))
let min_46360_73640 = minimum(v(n_46360_73640))
let min_46360_76440 = minimum(v(n_46360_76440))
let min_46360_79240 = minimum(v(n_46360_79240))
let min_46360_82040 = minimum(v(n_46360_82040))
let min_46360_84840 = minimum(v(n_46360_84840))
let min_46360_87640 = minimum(v(n_46360_87640))
let min_46740_40040 = minimum(v(n_46740_40040))
let min_46740_42840 = minimum(v(n_46740_42840))
let min_46740_45640 = minimum(v(n_46740_45640))
let min_46740_48440 = minimum(v(n_46740_48440))
let min_46740_51240 = minimum(v(n_46740_51240))
let min_46740_54040 = minimum(v(n_46740_54040))
let min_46740_56840 = minimum(v(n_46740_56840))
let min_46740_59640 = minimum(v(n_46740_59640))
let min_46740_62440 = minimum(v(n_46740_62440))
let min_46740_65240 = minimum(v(n_46740_65240))
let min_46740_68040 = minimum(v(n_46740_68040))
let min_46740_70840 = minimum(v(n_46740_70840))
let min_46740_73640 = minimum(v(n_46740_73640))
let min_46740_76440 = minimum(v(n_46740_76440))
let min_46740_79240 = minimum(v(n_46740_79240))
let min_46740_82040 = minimum(v(n_46740_82040))
let min_46740_84840 = minimum(v(n_46740_84840))
let min_46740_87640 = minimum(v(n_46740_87640))
let min_47120_40040 = minimum(v(n_47120_40040))
let min_47120_42840 = minimum(v(n_47120_42840))
let min_47120_45640 = minimum(v(n_47120_45640))
let min_47120_48440 = minimum(v(n_47120_48440))
let min_47120_51240 = minimum(v(n_47120_51240))
let min_47120_54040 = minimum(v(n_47120_54040))
let min_47120_56840 = minimum(v(n_47120_56840))
let min_47120_59640 = minimum(v(n_47120_59640))
let min_47120_62440 = minimum(v(n_47120_62440))
let min_47120_65240 = minimum(v(n_47120_65240))
let min_47120_68040 = minimum(v(n_47120_68040))
let min_47120_70840 = minimum(v(n_47120_70840))
let min_47120_73640 = minimum(v(n_47120_73640))
let min_47120_76440 = minimum(v(n_47120_76440))
let min_47120_79240 = minimum(v(n_47120_79240))
let min_47120_82040 = minimum(v(n_47120_82040))
let min_47120_84840 = minimum(v(n_47120_84840))
let min_47120_87640 = minimum(v(n_47120_87640))
let min_47500_40040 = minimum(v(n_47500_40040))
let min_47500_42840 = minimum(v(n_47500_42840))
let min_47500_45640 = minimum(v(n_47500_45640))
let min_47500_48440 = minimum(v(n_47500_48440))
let min_47500_51240 = minimum(v(n_47500_51240))
let min_47500_54040 = minimum(v(n_47500_54040))
let min_47500_56840 = minimum(v(n_47500_56840))
let min_47500_59640 = minimum(v(n_47500_59640))
let min_47500_62440 = minimum(v(n_47500_62440))
let min_47500_65240 = minimum(v(n_47500_65240))
let min_47500_68040 = minimum(v(n_47500_68040))
let min_47500_70840 = minimum(v(n_47500_70840))
let min_47500_73640 = minimum(v(n_47500_73640))
let min_47500_76440 = minimum(v(n_47500_76440))
let min_47500_79240 = minimum(v(n_47500_79240))
let min_47500_82040 = minimum(v(n_47500_82040))
let min_47500_84840 = minimum(v(n_47500_84840))
let min_47500_87640 = minimum(v(n_47500_87640))
let min_47880_40040 = minimum(v(n_47880_40040))
let min_47880_42840 = minimum(v(n_47880_42840))
let min_47880_45640 = minimum(v(n_47880_45640))
let min_47880_48440 = minimum(v(n_47880_48440))
let min_47880_51240 = minimum(v(n_47880_51240))
let min_47880_54040 = minimum(v(n_47880_54040))
let min_47880_56840 = minimum(v(n_47880_56840))
let min_47880_59640 = minimum(v(n_47880_59640))
let min_47880_62440 = minimum(v(n_47880_62440))
let min_47880_65240 = minimum(v(n_47880_65240))
let min_47880_68040 = minimum(v(n_47880_68040))
let min_47880_70840 = minimum(v(n_47880_70840))
let min_47880_73640 = minimum(v(n_47880_73640))
let min_47880_76440 = minimum(v(n_47880_76440))
let min_47880_79240 = minimum(v(n_47880_79240))
let min_47880_82040 = minimum(v(n_47880_82040))
let min_47880_84840 = minimum(v(n_47880_84840))
let min_47880_87640 = minimum(v(n_47880_87640))
let min_48260_40040 = minimum(v(n_48260_40040))
let min_48260_42840 = minimum(v(n_48260_42840))
let min_48260_45640 = minimum(v(n_48260_45640))
let min_48260_48440 = minimum(v(n_48260_48440))
let min_48260_51240 = minimum(v(n_48260_51240))
let min_48260_54040 = minimum(v(n_48260_54040))
let min_48260_56840 = minimum(v(n_48260_56840))
let min_48260_59640 = minimum(v(n_48260_59640))
let min_48260_62440 = minimum(v(n_48260_62440))
let min_48260_65240 = minimum(v(n_48260_65240))
let min_48260_68040 = minimum(v(n_48260_68040))
let min_48260_70840 = minimum(v(n_48260_70840))
let min_48260_73640 = minimum(v(n_48260_73640))
let min_48260_76440 = minimum(v(n_48260_76440))
let min_48260_79240 = minimum(v(n_48260_79240))
let min_48260_82040 = minimum(v(n_48260_82040))
let min_48260_84840 = minimum(v(n_48260_84840))
let min_48260_87640 = minimum(v(n_48260_87640))
let min_48640_40040 = minimum(v(n_48640_40040))
let min_48640_42840 = minimum(v(n_48640_42840))
let min_48640_45640 = minimum(v(n_48640_45640))
let min_48640_48440 = minimum(v(n_48640_48440))
let min_48640_51240 = minimum(v(n_48640_51240))
let min_48640_54040 = minimum(v(n_48640_54040))
let min_48640_56840 = minimum(v(n_48640_56840))
let min_48640_59640 = minimum(v(n_48640_59640))
let min_48640_62440 = minimum(v(n_48640_62440))
let min_48640_65240 = minimum(v(n_48640_65240))
let min_48640_68040 = minimum(v(n_48640_68040))
let min_48640_70840 = minimum(v(n_48640_70840))
let min_48640_73640 = minimum(v(n_48640_73640))
let min_48640_76440 = minimum(v(n_48640_76440))
let min_48640_79240 = minimum(v(n_48640_79240))
let min_48640_82040 = minimum(v(n_48640_82040))
let min_48640_84840 = minimum(v(n_48640_84840))
let min_48640_87640 = minimum(v(n_48640_87640))
let min_49020_40040 = minimum(v(n_49020_40040))
let min_49020_42840 = minimum(v(n_49020_42840))
let min_49020_45640 = minimum(v(n_49020_45640))
let min_49020_48440 = minimum(v(n_49020_48440))
let min_49020_51240 = minimum(v(n_49020_51240))
let min_49020_54040 = minimum(v(n_49020_54040))
let min_49020_56840 = minimum(v(n_49020_56840))
let min_49020_59640 = minimum(v(n_49020_59640))
let min_49020_62440 = minimum(v(n_49020_62440))
let min_49020_65240 = minimum(v(n_49020_65240))
let min_49020_68040 = minimum(v(n_49020_68040))
let min_49020_70840 = minimum(v(n_49020_70840))
let min_49020_73640 = minimum(v(n_49020_73640))
let min_49020_76440 = minimum(v(n_49020_76440))
let min_49020_79240 = minimum(v(n_49020_79240))
let min_49020_82040 = minimum(v(n_49020_82040))
let min_49020_84840 = minimum(v(n_49020_84840))
let min_49020_87640 = minimum(v(n_49020_87640))
let min_49400_40040 = minimum(v(n_49400_40040))
let min_49400_42840 = minimum(v(n_49400_42840))
let min_49400_45640 = minimum(v(n_49400_45640))
let min_49400_48440 = minimum(v(n_49400_48440))
let min_49400_51240 = minimum(v(n_49400_51240))
let min_49400_54040 = minimum(v(n_49400_54040))
let min_49400_56840 = minimum(v(n_49400_56840))
let min_49400_59640 = minimum(v(n_49400_59640))
let min_49400_62440 = minimum(v(n_49400_62440))
let min_49400_65240 = minimum(v(n_49400_65240))
let min_49400_68040 = minimum(v(n_49400_68040))
let min_49400_70840 = minimum(v(n_49400_70840))
let min_49400_73640 = minimum(v(n_49400_73640))
let min_49400_76440 = minimum(v(n_49400_76440))
let min_49400_79240 = minimum(v(n_49400_79240))
let min_49400_82040 = minimum(v(n_49400_82040))
let min_49400_84840 = minimum(v(n_49400_84840))
let min_49400_87640 = minimum(v(n_49400_87640))
let min_49780_40040 = minimum(v(n_49780_40040))
let min_49780_42840 = minimum(v(n_49780_42840))
let min_49780_45640 = minimum(v(n_49780_45640))
let min_49780_48440 = minimum(v(n_49780_48440))
let min_49780_51240 = minimum(v(n_49780_51240))
let min_49780_54040 = minimum(v(n_49780_54040))
let min_49780_56840 = minimum(v(n_49780_56840))
let min_49780_59640 = minimum(v(n_49780_59640))
let min_49780_62440 = minimum(v(n_49780_62440))
let min_49780_65240 = minimum(v(n_49780_65240))
let min_49780_68040 = minimum(v(n_49780_68040))
let min_49780_70840 = minimum(v(n_49780_70840))
let min_49780_73640 = minimum(v(n_49780_73640))
let min_49780_76440 = minimum(v(n_49780_76440))
let min_49780_79240 = minimum(v(n_49780_79240))
let min_49780_82040 = minimum(v(n_49780_82040))
let min_49780_84840 = minimum(v(n_49780_84840))
let min_49780_87640 = minimum(v(n_49780_87640))
let min_50160_40040 = minimum(v(n_50160_40040))
let min_50160_42840 = minimum(v(n_50160_42840))
let min_50160_45640 = minimum(v(n_50160_45640))
let min_50160_48440 = minimum(v(n_50160_48440))
let min_50160_51240 = minimum(v(n_50160_51240))
let min_50160_54040 = minimum(v(n_50160_54040))
let min_50160_56840 = minimum(v(n_50160_56840))
let min_50160_59640 = minimum(v(n_50160_59640))
let min_50160_62440 = minimum(v(n_50160_62440))
let min_50160_65240 = minimum(v(n_50160_65240))
let min_50160_68040 = minimum(v(n_50160_68040))
let min_50160_70840 = minimum(v(n_50160_70840))
let min_50160_73640 = minimum(v(n_50160_73640))
let min_50160_76440 = minimum(v(n_50160_76440))
let min_50160_79240 = minimum(v(n_50160_79240))
let min_50160_82040 = minimum(v(n_50160_82040))
let min_50160_84840 = minimum(v(n_50160_84840))
let min_50160_87640 = minimum(v(n_50160_87640))
let min_50540_40040 = minimum(v(n_50540_40040))
let min_50540_42840 = minimum(v(n_50540_42840))
let min_50540_45640 = minimum(v(n_50540_45640))
let min_50540_48440 = minimum(v(n_50540_48440))
let min_50540_51240 = minimum(v(n_50540_51240))
let min_50540_54040 = minimum(v(n_50540_54040))
let min_50540_56840 = minimum(v(n_50540_56840))
let min_50540_59640 = minimum(v(n_50540_59640))
let min_50540_62440 = minimum(v(n_50540_62440))
let min_50540_65240 = minimum(v(n_50540_65240))
let min_50540_68040 = minimum(v(n_50540_68040))
let min_50540_70840 = minimum(v(n_50540_70840))
let min_50540_73640 = minimum(v(n_50540_73640))
let min_50540_76440 = minimum(v(n_50540_76440))
let min_50540_79240 = minimum(v(n_50540_79240))
let min_50540_82040 = minimum(v(n_50540_82040))
let min_50540_84840 = minimum(v(n_50540_84840))
let min_50540_87640 = minimum(v(n_50540_87640))
let min_50920_40040 = minimum(v(n_50920_40040))
let min_50920_42840 = minimum(v(n_50920_42840))
let min_50920_45640 = minimum(v(n_50920_45640))
let min_50920_48440 = minimum(v(n_50920_48440))
let min_50920_51240 = minimum(v(n_50920_51240))
let min_50920_54040 = minimum(v(n_50920_54040))
let min_50920_56840 = minimum(v(n_50920_56840))
let min_50920_59640 = minimum(v(n_50920_59640))
let min_50920_62440 = minimum(v(n_50920_62440))
let min_50920_65240 = minimum(v(n_50920_65240))
let min_50920_68040 = minimum(v(n_50920_68040))
let min_50920_70840 = minimum(v(n_50920_70840))
let min_50920_73640 = minimum(v(n_50920_73640))
let min_50920_76440 = minimum(v(n_50920_76440))
let min_50920_79240 = minimum(v(n_50920_79240))
let min_50920_82040 = minimum(v(n_50920_82040))
let min_50920_84840 = minimum(v(n_50920_84840))
let min_50920_87640 = minimum(v(n_50920_87640))
let min_51300_40040 = minimum(v(n_51300_40040))
let min_51300_42840 = minimum(v(n_51300_42840))
let min_51300_45640 = minimum(v(n_51300_45640))
let min_51300_48440 = minimum(v(n_51300_48440))
let min_51300_51240 = minimum(v(n_51300_51240))
let min_51300_54040 = minimum(v(n_51300_54040))
let min_51300_56840 = minimum(v(n_51300_56840))
let min_51300_59640 = minimum(v(n_51300_59640))
let min_51300_62440 = minimum(v(n_51300_62440))
let min_51300_65240 = minimum(v(n_51300_65240))
let min_51300_68040 = minimum(v(n_51300_68040))
let min_51300_70840 = minimum(v(n_51300_70840))
let min_51300_73640 = minimum(v(n_51300_73640))
let min_51300_76440 = minimum(v(n_51300_76440))
let min_51300_79240 = minimum(v(n_51300_79240))
let min_51300_82040 = minimum(v(n_51300_82040))
let min_51300_84840 = minimum(v(n_51300_84840))
let min_51300_87640 = minimum(v(n_51300_87640))
let min_51680_40040 = minimum(v(n_51680_40040))
let min_51680_42840 = minimum(v(n_51680_42840))
let min_51680_45640 = minimum(v(n_51680_45640))
let min_51680_48440 = minimum(v(n_51680_48440))
let min_51680_51240 = minimum(v(n_51680_51240))
let min_51680_54040 = minimum(v(n_51680_54040))
let min_51680_56840 = minimum(v(n_51680_56840))
let min_51680_59640 = minimum(v(n_51680_59640))
let min_51680_62440 = minimum(v(n_51680_62440))
let min_51680_65240 = minimum(v(n_51680_65240))
let min_51680_68040 = minimum(v(n_51680_68040))
let min_51680_70840 = minimum(v(n_51680_70840))
let min_51680_73640 = minimum(v(n_51680_73640))
let min_51680_76440 = minimum(v(n_51680_76440))
let min_51680_79240 = minimum(v(n_51680_79240))
let min_51680_82040 = minimum(v(n_51680_82040))
let min_51680_84840 = minimum(v(n_51680_84840))
let min_51680_87640 = minimum(v(n_51680_87640))
let min_52060_40040 = minimum(v(n_52060_40040))
let min_52060_42840 = minimum(v(n_52060_42840))
let min_52060_45640 = minimum(v(n_52060_45640))
let min_52060_48440 = minimum(v(n_52060_48440))
let min_52060_51240 = minimum(v(n_52060_51240))
let min_52060_54040 = minimum(v(n_52060_54040))
let min_52060_56840 = minimum(v(n_52060_56840))
let min_52060_59640 = minimum(v(n_52060_59640))
let min_52060_62440 = minimum(v(n_52060_62440))
let min_52060_65240 = minimum(v(n_52060_65240))
let min_52060_68040 = minimum(v(n_52060_68040))
let min_52060_70840 = minimum(v(n_52060_70840))
let min_52060_73640 = minimum(v(n_52060_73640))
let min_52060_76440 = minimum(v(n_52060_76440))
let min_52060_79240 = minimum(v(n_52060_79240))
let min_52060_82040 = minimum(v(n_52060_82040))
let min_52060_84840 = minimum(v(n_52060_84840))
let min_52060_87640 = minimum(v(n_52060_87640))
let min_52440_40040 = minimum(v(n_52440_40040))
let min_52440_42840 = minimum(v(n_52440_42840))
let min_52440_45640 = minimum(v(n_52440_45640))
let min_52440_48440 = minimum(v(n_52440_48440))
let min_52440_51240 = minimum(v(n_52440_51240))
let min_52440_54040 = minimum(v(n_52440_54040))
let min_52440_56840 = minimum(v(n_52440_56840))
let min_52440_59640 = minimum(v(n_52440_59640))
let min_52440_62440 = minimum(v(n_52440_62440))
let min_52440_65240 = minimum(v(n_52440_65240))
let min_52440_68040 = minimum(v(n_52440_68040))
let min_52440_70840 = minimum(v(n_52440_70840))
let min_52440_73640 = minimum(v(n_52440_73640))
let min_52440_76440 = minimum(v(n_52440_76440))
let min_52440_79240 = minimum(v(n_52440_79240))
let min_52440_82040 = minimum(v(n_52440_82040))
let min_52440_84840 = minimum(v(n_52440_84840))
let min_52440_87640 = minimum(v(n_52440_87640))
let min_52820_40040 = minimum(v(n_52820_40040))
let min_52820_42840 = minimum(v(n_52820_42840))
let min_52820_45640 = minimum(v(n_52820_45640))
let min_52820_48440 = minimum(v(n_52820_48440))
let min_52820_51240 = minimum(v(n_52820_51240))
let min_52820_54040 = minimum(v(n_52820_54040))
let min_52820_56840 = minimum(v(n_52820_56840))
let min_52820_59640 = minimum(v(n_52820_59640))
let min_52820_62440 = minimum(v(n_52820_62440))
let min_52820_65240 = minimum(v(n_52820_65240))
let min_52820_68040 = minimum(v(n_52820_68040))
let min_52820_70840 = minimum(v(n_52820_70840))
let min_52820_73640 = minimum(v(n_52820_73640))
let min_52820_76440 = minimum(v(n_52820_76440))
let min_52820_79240 = minimum(v(n_52820_79240))
let min_52820_82040 = minimum(v(n_52820_82040))
let min_52820_84840 = minimum(v(n_52820_84840))
let min_52820_87640 = minimum(v(n_52820_87640))
let min_53200_40040 = minimum(v(n_53200_40040))
let min_53200_42840 = minimum(v(n_53200_42840))
let min_53200_45640 = minimum(v(n_53200_45640))
let min_53200_48440 = minimum(v(n_53200_48440))
let min_53200_51240 = minimum(v(n_53200_51240))
let min_53200_54040 = minimum(v(n_53200_54040))
let min_53200_56840 = minimum(v(n_53200_56840))
let min_53200_59640 = minimum(v(n_53200_59640))
let min_53200_62440 = minimum(v(n_53200_62440))
let min_53200_65240 = minimum(v(n_53200_65240))
let min_53200_68040 = minimum(v(n_53200_68040))
let min_53200_70840 = minimum(v(n_53200_70840))
let min_53200_73640 = minimum(v(n_53200_73640))
let min_53200_76440 = minimum(v(n_53200_76440))
let min_53200_79240 = minimum(v(n_53200_79240))
let min_53200_82040 = minimum(v(n_53200_82040))
let min_53200_84840 = minimum(v(n_53200_84840))
let min_53200_87640 = minimum(v(n_53200_87640))
let min_53580_40040 = minimum(v(n_53580_40040))
let min_53580_42840 = minimum(v(n_53580_42840))
let min_53580_45640 = minimum(v(n_53580_45640))
let min_53580_48440 = minimum(v(n_53580_48440))
let min_53580_51240 = minimum(v(n_53580_51240))
let min_53580_54040 = minimum(v(n_53580_54040))
let min_53580_56840 = minimum(v(n_53580_56840))
let min_53580_59640 = minimum(v(n_53580_59640))
let min_53580_62440 = minimum(v(n_53580_62440))
let min_53580_65240 = minimum(v(n_53580_65240))
let min_53580_68040 = minimum(v(n_53580_68040))
let min_53580_70840 = minimum(v(n_53580_70840))
let min_53580_73640 = minimum(v(n_53580_73640))
let min_53580_76440 = minimum(v(n_53580_76440))
let min_53580_79240 = minimum(v(n_53580_79240))
let min_53580_82040 = minimum(v(n_53580_82040))
let min_53580_84840 = minimum(v(n_53580_84840))
let min_53580_87640 = minimum(v(n_53580_87640))
let min_53960_40040 = minimum(v(n_53960_40040))
let min_53960_42840 = minimum(v(n_53960_42840))
let min_53960_45640 = minimum(v(n_53960_45640))
let min_53960_48440 = minimum(v(n_53960_48440))
let min_53960_51240 = minimum(v(n_53960_51240))
let min_53960_54040 = minimum(v(n_53960_54040))
let min_53960_56840 = minimum(v(n_53960_56840))
let min_53960_59640 = minimum(v(n_53960_59640))
let min_53960_62440 = minimum(v(n_53960_62440))
let min_53960_65240 = minimum(v(n_53960_65240))
let min_53960_68040 = minimum(v(n_53960_68040))
let min_53960_70840 = minimum(v(n_53960_70840))
let min_53960_73640 = minimum(v(n_53960_73640))
let min_53960_76440 = minimum(v(n_53960_76440))
let min_53960_79240 = minimum(v(n_53960_79240))
let min_53960_82040 = minimum(v(n_53960_82040))
let min_53960_84840 = minimum(v(n_53960_84840))
let min_53960_87640 = minimum(v(n_53960_87640))
let min_54340_40040 = minimum(v(n_54340_40040))
let min_54340_42840 = minimum(v(n_54340_42840))
let min_54340_45640 = minimum(v(n_54340_45640))
let min_54340_48440 = minimum(v(n_54340_48440))
let min_54340_51240 = minimum(v(n_54340_51240))
let min_54340_54040 = minimum(v(n_54340_54040))
let min_54340_56840 = minimum(v(n_54340_56840))
let min_54340_59640 = minimum(v(n_54340_59640))
let min_54340_62440 = minimum(v(n_54340_62440))
let min_54340_65240 = minimum(v(n_54340_65240))
let min_54340_68040 = minimum(v(n_54340_68040))
let min_54340_70840 = minimum(v(n_54340_70840))
let min_54340_73640 = minimum(v(n_54340_73640))
let min_54340_76440 = minimum(v(n_54340_76440))
let min_54340_79240 = minimum(v(n_54340_79240))
let min_54340_82040 = minimum(v(n_54340_82040))
let min_54340_84840 = minimum(v(n_54340_84840))
let min_54340_87640 = minimum(v(n_54340_87640))
let min_54720_40040 = minimum(v(n_54720_40040))
let min_54720_42840 = minimum(v(n_54720_42840))
let min_54720_45640 = minimum(v(n_54720_45640))
let min_54720_48440 = minimum(v(n_54720_48440))
let min_54720_51240 = minimum(v(n_54720_51240))
let min_54720_54040 = minimum(v(n_54720_54040))
let min_54720_56840 = minimum(v(n_54720_56840))
let min_54720_59640 = minimum(v(n_54720_59640))
let min_54720_62440 = minimum(v(n_54720_62440))
let min_54720_65240 = minimum(v(n_54720_65240))
let min_54720_68040 = minimum(v(n_54720_68040))
let min_54720_70840 = minimum(v(n_54720_70840))
let min_54720_73640 = minimum(v(n_54720_73640))
let min_54720_76440 = minimum(v(n_54720_76440))
let min_54720_79240 = minimum(v(n_54720_79240))
let min_54720_82040 = minimum(v(n_54720_82040))
let min_54720_84840 = minimum(v(n_54720_84840))
let min_54720_87640 = minimum(v(n_54720_87640))
let min_55100_40040 = minimum(v(n_55100_40040))
let min_55100_42840 = minimum(v(n_55100_42840))
let min_55100_45640 = minimum(v(n_55100_45640))
let min_55100_48440 = minimum(v(n_55100_48440))
let min_55100_51240 = minimum(v(n_55100_51240))
let min_55100_54040 = minimum(v(n_55100_54040))
let min_55100_56840 = minimum(v(n_55100_56840))
let min_55100_59640 = minimum(v(n_55100_59640))
let min_55100_62440 = minimum(v(n_55100_62440))
let min_55100_65240 = minimum(v(n_55100_65240))
let min_55100_68040 = minimum(v(n_55100_68040))
let min_55100_70840 = minimum(v(n_55100_70840))
let min_55100_73640 = minimum(v(n_55100_73640))
let min_55100_76440 = minimum(v(n_55100_76440))
let min_55100_79240 = minimum(v(n_55100_79240))
let min_55100_82040 = minimum(v(n_55100_82040))
let min_55100_84840 = minimum(v(n_55100_84840))
let min_55100_87640 = minimum(v(n_55100_87640))
let min_55480_40040 = minimum(v(n_55480_40040))
let min_55480_42840 = minimum(v(n_55480_42840))
let min_55480_45640 = minimum(v(n_55480_45640))
let min_55480_48440 = minimum(v(n_55480_48440))
let min_55480_51240 = minimum(v(n_55480_51240))
let min_55480_54040 = minimum(v(n_55480_54040))
let min_55480_56840 = minimum(v(n_55480_56840))
let min_55480_59640 = minimum(v(n_55480_59640))
let min_55480_62440 = minimum(v(n_55480_62440))
let min_55480_65240 = minimum(v(n_55480_65240))
let min_55480_68040 = minimum(v(n_55480_68040))
let min_55480_70840 = minimum(v(n_55480_70840))
let min_55480_73640 = minimum(v(n_55480_73640))
let min_55480_76440 = minimum(v(n_55480_76440))
let min_55480_79240 = minimum(v(n_55480_79240))
let min_55480_82040 = minimum(v(n_55480_82040))
let min_55480_84840 = minimum(v(n_55480_84840))
let min_55480_87640 = minimum(v(n_55480_87640))
let min_55860_40040 = minimum(v(n_55860_40040))
let min_55860_42840 = minimum(v(n_55860_42840))
let min_55860_45640 = minimum(v(n_55860_45640))
let min_55860_48440 = minimum(v(n_55860_48440))
let min_55860_51240 = minimum(v(n_55860_51240))
let min_55860_54040 = minimum(v(n_55860_54040))
let min_55860_56840 = minimum(v(n_55860_56840))
let min_55860_59640 = minimum(v(n_55860_59640))
let min_55860_62440 = minimum(v(n_55860_62440))
let min_55860_65240 = minimum(v(n_55860_65240))
let min_55860_68040 = minimum(v(n_55860_68040))
let min_55860_70840 = minimum(v(n_55860_70840))
let min_55860_73640 = minimum(v(n_55860_73640))
let min_55860_76440 = minimum(v(n_55860_76440))
let min_55860_79240 = minimum(v(n_55860_79240))
let min_55860_82040 = minimum(v(n_55860_82040))
let min_55860_84840 = minimum(v(n_55860_84840))
let min_55860_87640 = minimum(v(n_55860_87640))
let min_56240_40040 = minimum(v(n_56240_40040))
let min_56240_42840 = minimum(v(n_56240_42840))
let min_56240_45640 = minimum(v(n_56240_45640))
let min_56240_48440 = minimum(v(n_56240_48440))
let min_56240_51240 = minimum(v(n_56240_51240))
let min_56240_54040 = minimum(v(n_56240_54040))
let min_56240_56840 = minimum(v(n_56240_56840))
let min_56240_59640 = minimum(v(n_56240_59640))
let min_56240_62440 = minimum(v(n_56240_62440))
let min_56240_65240 = minimum(v(n_56240_65240))
let min_56240_68040 = minimum(v(n_56240_68040))
let min_56240_70840 = minimum(v(n_56240_70840))
let min_56240_73640 = minimum(v(n_56240_73640))
let min_56240_76440 = minimum(v(n_56240_76440))
let min_56240_79240 = minimum(v(n_56240_79240))
let min_56240_82040 = minimum(v(n_56240_82040))
let min_56240_84840 = minimum(v(n_56240_84840))
let min_56240_87640 = minimum(v(n_56240_87640))
let min_56620_40040 = minimum(v(n_56620_40040))
let min_56620_42840 = minimum(v(n_56620_42840))
let min_56620_45640 = minimum(v(n_56620_45640))
let min_56620_48440 = minimum(v(n_56620_48440))
let min_56620_51240 = minimum(v(n_56620_51240))
let min_56620_54040 = minimum(v(n_56620_54040))
let min_56620_56840 = minimum(v(n_56620_56840))
let min_56620_59640 = minimum(v(n_56620_59640))
let min_56620_62440 = minimum(v(n_56620_62440))
let min_56620_65240 = minimum(v(n_56620_65240))
let min_56620_68040 = minimum(v(n_56620_68040))
let min_56620_70840 = minimum(v(n_56620_70840))
let min_56620_73640 = minimum(v(n_56620_73640))
let min_56620_76440 = minimum(v(n_56620_76440))
let min_56620_79240 = minimum(v(n_56620_79240))
let min_56620_82040 = minimum(v(n_56620_82040))
let min_56620_84840 = minimum(v(n_56620_84840))
let min_56620_87640 = minimum(v(n_56620_87640))
let min_57000_40040 = minimum(v(n_57000_40040))
let min_57000_42840 = minimum(v(n_57000_42840))
let min_57000_45640 = minimum(v(n_57000_45640))
let min_57000_48440 = minimum(v(n_57000_48440))
let min_57000_51240 = minimum(v(n_57000_51240))
let min_57000_54040 = minimum(v(n_57000_54040))
let min_57000_56840 = minimum(v(n_57000_56840))
let min_57000_59640 = minimum(v(n_57000_59640))
let min_57000_62440 = minimum(v(n_57000_62440))
let min_57000_65240 = minimum(v(n_57000_65240))
let min_57000_68040 = minimum(v(n_57000_68040))
let min_57000_70840 = minimum(v(n_57000_70840))
let min_57000_73640 = minimum(v(n_57000_73640))
let min_57000_76440 = minimum(v(n_57000_76440))
let min_57000_79240 = minimum(v(n_57000_79240))
let min_57000_82040 = minimum(v(n_57000_82040))
let min_57000_84840 = minimum(v(n_57000_84840))
let min_57000_87640 = minimum(v(n_57000_87640))
let min_57380_40040 = minimum(v(n_57380_40040))
let min_57380_42840 = minimum(v(n_57380_42840))
let min_57380_45640 = minimum(v(n_57380_45640))
let min_57380_48440 = minimum(v(n_57380_48440))
let min_57380_51240 = minimum(v(n_57380_51240))
let min_57380_54040 = minimum(v(n_57380_54040))
let min_57380_56840 = minimum(v(n_57380_56840))
let min_57380_59640 = minimum(v(n_57380_59640))
let min_57380_62440 = minimum(v(n_57380_62440))
let min_57380_65240 = minimum(v(n_57380_65240))
let min_57380_68040 = minimum(v(n_57380_68040))
let min_57380_70840 = minimum(v(n_57380_70840))
let min_57380_73640 = minimum(v(n_57380_73640))
let min_57380_76440 = minimum(v(n_57380_76440))
let min_57380_79240 = minimum(v(n_57380_79240))
let min_57380_82040 = minimum(v(n_57380_82040))
let min_57380_84840 = minimum(v(n_57380_84840))
let min_57380_87640 = minimum(v(n_57380_87640))
let min_57760_40040 = minimum(v(n_57760_40040))
let min_57760_42840 = minimum(v(n_57760_42840))
let min_57760_45640 = minimum(v(n_57760_45640))
let min_57760_48440 = minimum(v(n_57760_48440))
let min_57760_51240 = minimum(v(n_57760_51240))
let min_57760_54040 = minimum(v(n_57760_54040))
let min_57760_56840 = minimum(v(n_57760_56840))
let min_57760_59640 = minimum(v(n_57760_59640))
let min_57760_62440 = minimum(v(n_57760_62440))
let min_57760_65240 = minimum(v(n_57760_65240))
let min_57760_68040 = minimum(v(n_57760_68040))
let min_57760_70840 = minimum(v(n_57760_70840))
let min_57760_73640 = minimum(v(n_57760_73640))
let min_57760_76440 = minimum(v(n_57760_76440))
let min_57760_79240 = minimum(v(n_57760_79240))
let min_57760_82040 = minimum(v(n_57760_82040))
let min_57760_84840 = minimum(v(n_57760_84840))
let min_57760_87640 = minimum(v(n_57760_87640))
let min_58140_40040 = minimum(v(n_58140_40040))
let min_58140_42840 = minimum(v(n_58140_42840))
let min_58140_45640 = minimum(v(n_58140_45640))
let min_58140_48440 = minimum(v(n_58140_48440))
let min_58140_51240 = minimum(v(n_58140_51240))
let min_58140_54040 = minimum(v(n_58140_54040))
let min_58140_56840 = minimum(v(n_58140_56840))
let min_58140_59640 = minimum(v(n_58140_59640))
let min_58140_62440 = minimum(v(n_58140_62440))
let min_58140_65240 = minimum(v(n_58140_65240))
let min_58140_68040 = minimum(v(n_58140_68040))
let min_58140_70840 = minimum(v(n_58140_70840))
let min_58140_73640 = minimum(v(n_58140_73640))
let min_58140_76440 = minimum(v(n_58140_76440))
let min_58140_79240 = minimum(v(n_58140_79240))
let min_58140_82040 = minimum(v(n_58140_82040))
let min_58140_84840 = minimum(v(n_58140_84840))
let min_58140_87640 = minimum(v(n_58140_87640))
let min_58520_40040 = minimum(v(n_58520_40040))
let min_58520_42840 = minimum(v(n_58520_42840))
let min_58520_45640 = minimum(v(n_58520_45640))
let min_58520_48440 = minimum(v(n_58520_48440))
let min_58520_51240 = minimum(v(n_58520_51240))
let min_58520_54040 = minimum(v(n_58520_54040))
let min_58520_56840 = minimum(v(n_58520_56840))
let min_58520_59640 = minimum(v(n_58520_59640))
let min_58520_62440 = minimum(v(n_58520_62440))
let min_58520_65240 = minimum(v(n_58520_65240))
let min_58520_68040 = minimum(v(n_58520_68040))
let min_58520_70840 = minimum(v(n_58520_70840))
let min_58520_73640 = minimum(v(n_58520_73640))
let min_58520_76440 = minimum(v(n_58520_76440))
let min_58520_79240 = minimum(v(n_58520_79240))
let min_58520_82040 = minimum(v(n_58520_82040))
let min_58520_84840 = minimum(v(n_58520_84840))
let min_58520_87640 = minimum(v(n_58520_87640))
let min_58900_40040 = minimum(v(n_58900_40040))
let min_58900_42840 = minimum(v(n_58900_42840))
let min_58900_45640 = minimum(v(n_58900_45640))
let min_58900_48440 = minimum(v(n_58900_48440))
let min_58900_51240 = minimum(v(n_58900_51240))
let min_58900_54040 = minimum(v(n_58900_54040))
let min_58900_56840 = minimum(v(n_58900_56840))
let min_58900_59640 = minimum(v(n_58900_59640))
let min_58900_62440 = minimum(v(n_58900_62440))
let min_58900_65240 = minimum(v(n_58900_65240))
let min_58900_68040 = minimum(v(n_58900_68040))
let min_58900_70840 = minimum(v(n_58900_70840))
let min_58900_73640 = minimum(v(n_58900_73640))
let min_58900_76440 = minimum(v(n_58900_76440))
let min_58900_79240 = minimum(v(n_58900_79240))
let min_58900_82040 = minimum(v(n_58900_82040))
let min_58900_84840 = minimum(v(n_58900_84840))
let min_58900_87640 = minimum(v(n_58900_87640))
let min_59280_40040 = minimum(v(n_59280_40040))
let min_59280_42840 = minimum(v(n_59280_42840))
let min_59280_45640 = minimum(v(n_59280_45640))
let min_59280_48440 = minimum(v(n_59280_48440))
let min_59280_51240 = minimum(v(n_59280_51240))
let min_59280_54040 = minimum(v(n_59280_54040))
let min_59280_56840 = minimum(v(n_59280_56840))
let min_59280_59640 = minimum(v(n_59280_59640))
let min_59280_62440 = minimum(v(n_59280_62440))
let min_59280_65240 = minimum(v(n_59280_65240))
let min_59280_68040 = minimum(v(n_59280_68040))
let min_59280_70840 = minimum(v(n_59280_70840))
let min_59280_73640 = minimum(v(n_59280_73640))
let min_59280_76440 = minimum(v(n_59280_76440))
let min_59280_79240 = minimum(v(n_59280_79240))
let min_59280_82040 = minimum(v(n_59280_82040))
let min_59280_84840 = minimum(v(n_59280_84840))
let min_59280_87640 = minimum(v(n_59280_87640))
let min_59660_40040 = minimum(v(n_59660_40040))
let min_59660_42840 = minimum(v(n_59660_42840))
let min_59660_45640 = minimum(v(n_59660_45640))
let min_59660_48440 = minimum(v(n_59660_48440))
let min_59660_51240 = minimum(v(n_59660_51240))
let min_59660_54040 = minimum(v(n_59660_54040))
let min_59660_56840 = minimum(v(n_59660_56840))
let min_59660_59640 = minimum(v(n_59660_59640))
let min_59660_62440 = minimum(v(n_59660_62440))
let min_59660_65240 = minimum(v(n_59660_65240))
let min_59660_68040 = minimum(v(n_59660_68040))
let min_59660_70840 = minimum(v(n_59660_70840))
let min_59660_73640 = minimum(v(n_59660_73640))
let min_59660_76440 = minimum(v(n_59660_76440))
let min_59660_79240 = minimum(v(n_59660_79240))
let min_59660_82040 = minimum(v(n_59660_82040))
let min_59660_84840 = minimum(v(n_59660_84840))
let min_59660_87640 = minimum(v(n_59660_87640))
let min_60040_40040 = minimum(v(n_60040_40040))
let min_60040_42840 = minimum(v(n_60040_42840))
let min_60040_45640 = minimum(v(n_60040_45640))
let min_60040_48440 = minimum(v(n_60040_48440))
let min_60040_51240 = minimum(v(n_60040_51240))
let min_60040_54040 = minimum(v(n_60040_54040))
let min_60040_56840 = minimum(v(n_60040_56840))
let min_60040_59640 = minimum(v(n_60040_59640))
let min_60040_62440 = minimum(v(n_60040_62440))
let min_60040_65240 = minimum(v(n_60040_65240))
let min_60040_68040 = minimum(v(n_60040_68040))
let min_60040_70840 = minimum(v(n_60040_70840))
let min_60040_73640 = minimum(v(n_60040_73640))
let min_60040_76440 = minimum(v(n_60040_76440))
let min_60040_79240 = minimum(v(n_60040_79240))
let min_60040_82040 = minimum(v(n_60040_82040))
let min_60040_84840 = minimum(v(n_60040_84840))
let min_60040_87640 = minimum(v(n_60040_87640))
let min_60420_40040 = minimum(v(n_60420_40040))
let min_60420_42840 = minimum(v(n_60420_42840))
let min_60420_45640 = minimum(v(n_60420_45640))
let min_60420_48440 = minimum(v(n_60420_48440))
let min_60420_51240 = minimum(v(n_60420_51240))
let min_60420_54040 = minimum(v(n_60420_54040))
let min_60420_56840 = minimum(v(n_60420_56840))
let min_60420_59640 = minimum(v(n_60420_59640))
let min_60420_62440 = minimum(v(n_60420_62440))
let min_60420_65240 = minimum(v(n_60420_65240))
let min_60420_68040 = minimum(v(n_60420_68040))
let min_60420_70840 = minimum(v(n_60420_70840))
let min_60420_73640 = minimum(v(n_60420_73640))
let min_60420_76440 = minimum(v(n_60420_76440))
let min_60420_79240 = minimum(v(n_60420_79240))
let min_60420_82040 = minimum(v(n_60420_82040))
let min_60420_84840 = minimum(v(n_60420_84840))
let min_60420_87640 = minimum(v(n_60420_87640))
let min_60800_40040 = minimum(v(n_60800_40040))
let min_60800_42840 = minimum(v(n_60800_42840))
let min_60800_45640 = minimum(v(n_60800_45640))
let min_60800_48440 = minimum(v(n_60800_48440))
let min_60800_51240 = minimum(v(n_60800_51240))
let min_60800_54040 = minimum(v(n_60800_54040))
let min_60800_56840 = minimum(v(n_60800_56840))
let min_60800_59640 = minimum(v(n_60800_59640))
let min_60800_62440 = minimum(v(n_60800_62440))
let min_60800_65240 = minimum(v(n_60800_65240))
let min_60800_68040 = minimum(v(n_60800_68040))
let min_60800_70840 = minimum(v(n_60800_70840))
let min_60800_73640 = minimum(v(n_60800_73640))
let min_60800_76440 = minimum(v(n_60800_76440))
let min_60800_79240 = minimum(v(n_60800_79240))
let min_60800_82040 = minimum(v(n_60800_82040))
let min_60800_84840 = minimum(v(n_60800_84840))
let min_60800_87640 = minimum(v(n_60800_87640))
let min_61180_40040 = minimum(v(n_61180_40040))
let min_61180_42840 = minimum(v(n_61180_42840))
let min_61180_45640 = minimum(v(n_61180_45640))
let min_61180_48440 = minimum(v(n_61180_48440))
let min_61180_51240 = minimum(v(n_61180_51240))
let min_61180_54040 = minimum(v(n_61180_54040))
let min_61180_56840 = minimum(v(n_61180_56840))
let min_61180_59640 = minimum(v(n_61180_59640))
let min_61180_62440 = minimum(v(n_61180_62440))
let min_61180_65240 = minimum(v(n_61180_65240))
let min_61180_68040 = minimum(v(n_61180_68040))
let min_61180_70840 = minimum(v(n_61180_70840))
let min_61180_73640 = minimum(v(n_61180_73640))
let min_61180_76440 = minimum(v(n_61180_76440))
let min_61180_79240 = minimum(v(n_61180_79240))
let min_61180_82040 = minimum(v(n_61180_82040))
let min_61180_84840 = minimum(v(n_61180_84840))
let min_61180_87640 = minimum(v(n_61180_87640))
let min_61560_40040 = minimum(v(n_61560_40040))
let min_61560_42840 = minimum(v(n_61560_42840))
let min_61560_45640 = minimum(v(n_61560_45640))
let min_61560_48440 = minimum(v(n_61560_48440))
let min_61560_51240 = minimum(v(n_61560_51240))
let min_61560_54040 = minimum(v(n_61560_54040))
let min_61560_56840 = minimum(v(n_61560_56840))
let min_61560_59640 = minimum(v(n_61560_59640))
let min_61560_62440 = minimum(v(n_61560_62440))
let min_61560_65240 = minimum(v(n_61560_65240))
let min_61560_68040 = minimum(v(n_61560_68040))
let min_61560_70840 = minimum(v(n_61560_70840))
let min_61560_73640 = minimum(v(n_61560_73640))
let min_61560_76440 = minimum(v(n_61560_76440))
let min_61560_79240 = minimum(v(n_61560_79240))
let min_61560_82040 = minimum(v(n_61560_82040))
let min_61560_84840 = minimum(v(n_61560_84840))
let min_61560_87640 = minimum(v(n_61560_87640))
let min_61940_40040 = minimum(v(n_61940_40040))
let min_61940_42840 = minimum(v(n_61940_42840))
let min_61940_45640 = minimum(v(n_61940_45640))
let min_61940_48440 = minimum(v(n_61940_48440))
let min_61940_51240 = minimum(v(n_61940_51240))
let min_61940_54040 = minimum(v(n_61940_54040))
let min_61940_56840 = minimum(v(n_61940_56840))
let min_61940_59640 = minimum(v(n_61940_59640))
let min_61940_62440 = minimum(v(n_61940_62440))
let min_61940_65240 = minimum(v(n_61940_65240))
let min_61940_68040 = minimum(v(n_61940_68040))
let min_61940_70840 = minimum(v(n_61940_70840))
let min_61940_73640 = minimum(v(n_61940_73640))
let min_61940_76440 = minimum(v(n_61940_76440))
let min_61940_79240 = minimum(v(n_61940_79240))
let min_61940_82040 = minimum(v(n_61940_82040))
let min_61940_84840 = minimum(v(n_61940_84840))
let min_61940_87640 = minimum(v(n_61940_87640))
let min_62320_40040 = minimum(v(n_62320_40040))
let min_62320_42840 = minimum(v(n_62320_42840))
let min_62320_45640 = minimum(v(n_62320_45640))
let min_62320_48440 = minimum(v(n_62320_48440))
let min_62320_51240 = minimum(v(n_62320_51240))
let min_62320_54040 = minimum(v(n_62320_54040))
let min_62320_56840 = minimum(v(n_62320_56840))
let min_62320_59640 = minimum(v(n_62320_59640))
let min_62320_62440 = minimum(v(n_62320_62440))
let min_62320_65240 = minimum(v(n_62320_65240))
let min_62320_68040 = minimum(v(n_62320_68040))
let min_62320_70840 = minimum(v(n_62320_70840))
let min_62320_73640 = minimum(v(n_62320_73640))
let min_62320_76440 = minimum(v(n_62320_76440))
let min_62320_79240 = minimum(v(n_62320_79240))
let min_62320_82040 = minimum(v(n_62320_82040))
let min_62320_84840 = minimum(v(n_62320_84840))
let min_62320_87640 = minimum(v(n_62320_87640))
let min_63080_40040 = minimum(v(n_63080_40040))
let min_63080_42840 = minimum(v(n_63080_42840))
let min_63080_45640 = minimum(v(n_63080_45640))
let min_63080_48440 = minimum(v(n_63080_48440))
let min_63080_51240 = minimum(v(n_63080_51240))
let min_63080_54040 = minimum(v(n_63080_54040))
let min_63080_56840 = minimum(v(n_63080_56840))
let min_63080_59640 = minimum(v(n_63080_59640))
let min_63080_62440 = minimum(v(n_63080_62440))
let min_63080_65240 = minimum(v(n_63080_65240))
let min_63080_68040 = minimum(v(n_63080_68040))
let min_63080_70840 = minimum(v(n_63080_70840))
let min_63080_73640 = minimum(v(n_63080_73640))
let min_63080_76440 = minimum(v(n_63080_76440))
let min_63080_79240 = minimum(v(n_63080_79240))
let min_63080_82040 = minimum(v(n_63080_82040))
let min_63080_84840 = minimum(v(n_63080_84840))
let min_63080_87640 = minimum(v(n_63080_87640))
let min_63460_40040 = minimum(v(n_63460_40040))
let min_63460_42840 = minimum(v(n_63460_42840))
let min_63460_45640 = minimum(v(n_63460_45640))
let min_63460_48440 = minimum(v(n_63460_48440))
let min_63460_51240 = minimum(v(n_63460_51240))
let min_63460_54040 = minimum(v(n_63460_54040))
let min_63460_56840 = minimum(v(n_63460_56840))
let min_63460_59640 = minimum(v(n_63460_59640))
let min_63460_62440 = minimum(v(n_63460_62440))
let min_63460_65240 = minimum(v(n_63460_65240))
let min_63460_68040 = minimum(v(n_63460_68040))
let min_63460_70840 = minimum(v(n_63460_70840))
let min_63460_73640 = minimum(v(n_63460_73640))
let min_63460_76440 = minimum(v(n_63460_76440))
let min_63460_79240 = minimum(v(n_63460_79240))
let min_63460_82040 = minimum(v(n_63460_82040))
let min_63460_84840 = minimum(v(n_63460_84840))
let min_63460_87640 = minimum(v(n_63460_87640))
let min_63840_40040 = minimum(v(n_63840_40040))
let min_63840_42840 = minimum(v(n_63840_42840))
let min_63840_45640 = minimum(v(n_63840_45640))
let min_63840_48440 = minimum(v(n_63840_48440))
let min_63840_51240 = minimum(v(n_63840_51240))
let min_63840_54040 = minimum(v(n_63840_54040))
let min_63840_56840 = minimum(v(n_63840_56840))
let min_63840_59640 = minimum(v(n_63840_59640))
let min_63840_62440 = minimum(v(n_63840_62440))
let min_63840_65240 = minimum(v(n_63840_65240))
let min_63840_68040 = minimum(v(n_63840_68040))
let min_63840_70840 = minimum(v(n_63840_70840))
let min_63840_73640 = minimum(v(n_63840_73640))
let min_63840_76440 = minimum(v(n_63840_76440))
let min_63840_79240 = minimum(v(n_63840_79240))
let min_63840_82040 = minimum(v(n_63840_82040))
let min_63840_84840 = minimum(v(n_63840_84840))
let min_63840_87640 = minimum(v(n_63840_87640))
let min_64220_40040 = minimum(v(n_64220_40040))
let min_64220_42840 = minimum(v(n_64220_42840))
let min_64220_45640 = minimum(v(n_64220_45640))
let min_64220_48440 = minimum(v(n_64220_48440))
let min_64220_51240 = minimum(v(n_64220_51240))
let min_64220_54040 = minimum(v(n_64220_54040))
let min_64220_56840 = minimum(v(n_64220_56840))
let min_64220_59640 = minimum(v(n_64220_59640))
let min_64220_62440 = minimum(v(n_64220_62440))
let min_64220_65240 = minimum(v(n_64220_65240))
let min_64220_68040 = minimum(v(n_64220_68040))
let min_64220_70840 = minimum(v(n_64220_70840))
let min_64220_73640 = minimum(v(n_64220_73640))
let min_64220_76440 = minimum(v(n_64220_76440))
let min_64220_79240 = minimum(v(n_64220_79240))
let min_64220_82040 = minimum(v(n_64220_82040))
let min_64220_84840 = minimum(v(n_64220_84840))
let min_64220_87640 = minimum(v(n_64220_87640))
let min_64600_40040 = minimum(v(n_64600_40040))
let min_64600_42840 = minimum(v(n_64600_42840))
let min_64600_45640 = minimum(v(n_64600_45640))
let min_64600_48440 = minimum(v(n_64600_48440))
let min_64600_51240 = minimum(v(n_64600_51240))
let min_64600_54040 = minimum(v(n_64600_54040))
let min_64600_56840 = minimum(v(n_64600_56840))
let min_64600_59640 = minimum(v(n_64600_59640))
let min_64600_62440 = minimum(v(n_64600_62440))
let min_64600_65240 = minimum(v(n_64600_65240))
let min_64600_68040 = minimum(v(n_64600_68040))
let min_64600_70840 = minimum(v(n_64600_70840))
let min_64600_73640 = minimum(v(n_64600_73640))
let min_64600_76440 = minimum(v(n_64600_76440))
let min_64600_79240 = minimum(v(n_64600_79240))
let min_64600_82040 = minimum(v(n_64600_82040))
let min_64600_84840 = minimum(v(n_64600_84840))
let min_64600_87640 = minimum(v(n_64600_87640))
let min_64980_40040 = minimum(v(n_64980_40040))
let min_64980_42840 = minimum(v(n_64980_42840))
let min_64980_45640 = minimum(v(n_64980_45640))
let min_64980_48440 = minimum(v(n_64980_48440))
let min_64980_51240 = minimum(v(n_64980_51240))
let min_64980_54040 = minimum(v(n_64980_54040))
let min_64980_56840 = minimum(v(n_64980_56840))
let min_64980_59640 = minimum(v(n_64980_59640))
let min_64980_62440 = minimum(v(n_64980_62440))
let min_64980_65240 = minimum(v(n_64980_65240))
let min_64980_68040 = minimum(v(n_64980_68040))
let min_64980_70840 = minimum(v(n_64980_70840))
let min_64980_73640 = minimum(v(n_64980_73640))
let min_64980_76440 = minimum(v(n_64980_76440))
let min_64980_79240 = minimum(v(n_64980_79240))
let min_64980_82040 = minimum(v(n_64980_82040))
let min_64980_84840 = minimum(v(n_64980_84840))
let min_64980_87640 = minimum(v(n_64980_87640))
let min_65360_40040 = minimum(v(n_65360_40040))
let min_65360_42840 = minimum(v(n_65360_42840))
let min_65360_45640 = minimum(v(n_65360_45640))
let min_65360_48440 = minimum(v(n_65360_48440))
let min_65360_51240 = minimum(v(n_65360_51240))
let min_65360_54040 = minimum(v(n_65360_54040))
let min_65360_56840 = minimum(v(n_65360_56840))
let min_65360_59640 = minimum(v(n_65360_59640))
let min_65360_62440 = minimum(v(n_65360_62440))
let min_65360_65240 = minimum(v(n_65360_65240))
let min_65360_68040 = minimum(v(n_65360_68040))
let min_65360_70840 = minimum(v(n_65360_70840))
let min_65360_73640 = minimum(v(n_65360_73640))
let min_65360_76440 = minimum(v(n_65360_76440))
let min_65360_79240 = minimum(v(n_65360_79240))
let min_65360_82040 = minimum(v(n_65360_82040))
let min_65360_84840 = minimum(v(n_65360_84840))
let min_65360_87640 = minimum(v(n_65360_87640))
let min_65740_40040 = minimum(v(n_65740_40040))
let min_65740_42840 = minimum(v(n_65740_42840))
let min_65740_45640 = minimum(v(n_65740_45640))
let min_65740_48440 = minimum(v(n_65740_48440))
let min_65740_51240 = minimum(v(n_65740_51240))
let min_65740_54040 = minimum(v(n_65740_54040))
let min_65740_56840 = minimum(v(n_65740_56840))
let min_65740_59640 = minimum(v(n_65740_59640))
let min_65740_62440 = minimum(v(n_65740_62440))
let min_65740_65240 = minimum(v(n_65740_65240))
let min_65740_68040 = minimum(v(n_65740_68040))
let min_65740_70840 = minimum(v(n_65740_70840))
let min_65740_73640 = minimum(v(n_65740_73640))
let min_65740_76440 = minimum(v(n_65740_76440))
let min_65740_79240 = minimum(v(n_65740_79240))
let min_65740_82040 = minimum(v(n_65740_82040))
let min_65740_84840 = minimum(v(n_65740_84840))
let min_65740_87640 = minimum(v(n_65740_87640))
let min_66120_40040 = minimum(v(n_66120_40040))
let min_66120_42840 = minimum(v(n_66120_42840))
let min_66120_45640 = minimum(v(n_66120_45640))
let min_66120_48440 = minimum(v(n_66120_48440))
let min_66120_51240 = minimum(v(n_66120_51240))
let min_66120_54040 = minimum(v(n_66120_54040))
let min_66120_56840 = minimum(v(n_66120_56840))
let min_66120_59640 = minimum(v(n_66120_59640))
let min_66120_62440 = minimum(v(n_66120_62440))
let min_66120_65240 = minimum(v(n_66120_65240))
let min_66120_68040 = minimum(v(n_66120_68040))
let min_66120_70840 = minimum(v(n_66120_70840))
let min_66120_73640 = minimum(v(n_66120_73640))
let min_66120_76440 = minimum(v(n_66120_76440))
let min_66120_79240 = minimum(v(n_66120_79240))
let min_66120_82040 = minimum(v(n_66120_82040))
let min_66120_84840 = minimum(v(n_66120_84840))
let min_66120_87640 = minimum(v(n_66120_87640))
let min_66880_40040 = minimum(v(n_66880_40040))
let min_66880_42840 = minimum(v(n_66880_42840))
let min_66880_45640 = minimum(v(n_66880_45640))
let min_66880_48440 = minimum(v(n_66880_48440))
let min_66880_51240 = minimum(v(n_66880_51240))
let min_66880_54040 = minimum(v(n_66880_54040))
let min_66880_56840 = minimum(v(n_66880_56840))
let min_66880_59640 = minimum(v(n_66880_59640))
let min_66880_62440 = minimum(v(n_66880_62440))
let min_66880_65240 = minimum(v(n_66880_65240))
let min_66880_68040 = minimum(v(n_66880_68040))
let min_66880_70840 = minimum(v(n_66880_70840))
let min_66880_73640 = minimum(v(n_66880_73640))
let min_66880_76440 = minimum(v(n_66880_76440))
let min_66880_79240 = minimum(v(n_66880_79240))
let min_66880_82040 = minimum(v(n_66880_82040))
let min_66880_84840 = minimum(v(n_66880_84840))
let min_66880_87640 = minimum(v(n_66880_87640))
let min_67260_40040 = minimum(v(n_67260_40040))
let min_67260_42840 = minimum(v(n_67260_42840))
let min_67260_45640 = minimum(v(n_67260_45640))
let min_67260_48440 = minimum(v(n_67260_48440))
let min_67260_51240 = minimum(v(n_67260_51240))
let min_67260_54040 = minimum(v(n_67260_54040))
let min_67260_56840 = minimum(v(n_67260_56840))
let min_67260_59640 = minimum(v(n_67260_59640))
let min_67260_62440 = minimum(v(n_67260_62440))
let min_67260_65240 = minimum(v(n_67260_65240))
let min_67260_68040 = minimum(v(n_67260_68040))
let min_67260_70840 = minimum(v(n_67260_70840))
let min_67260_73640 = minimum(v(n_67260_73640))
let min_67260_76440 = minimum(v(n_67260_76440))
let min_67260_79240 = minimum(v(n_67260_79240))
let min_67260_82040 = minimum(v(n_67260_82040))
let min_67260_84840 = minimum(v(n_67260_84840))
let min_67260_87640 = minimum(v(n_67260_87640))
let min_68020_40040 = minimum(v(n_68020_40040))
let min_68020_42840 = minimum(v(n_68020_42840))
let min_68020_45640 = minimum(v(n_68020_45640))
let min_68020_48440 = minimum(v(n_68020_48440))
let min_68020_51240 = minimum(v(n_68020_51240))
let min_68020_54040 = minimum(v(n_68020_54040))
let min_68020_56840 = minimum(v(n_68020_56840))
let min_68020_59640 = minimum(v(n_68020_59640))
let min_68020_62440 = minimum(v(n_68020_62440))
let min_68020_65240 = minimum(v(n_68020_65240))
let min_68020_68040 = minimum(v(n_68020_68040))
let min_68020_70840 = minimum(v(n_68020_70840))
let min_68020_73640 = minimum(v(n_68020_73640))
let min_68020_76440 = minimum(v(n_68020_76440))
let min_68020_79240 = minimum(v(n_68020_79240))
let min_68020_82040 = minimum(v(n_68020_82040))
let min_68020_84840 = minimum(v(n_68020_84840))
let min_68020_87640 = minimum(v(n_68020_87640))
let min_68400_40040 = minimum(v(n_68400_40040))
let min_68400_42840 = minimum(v(n_68400_42840))
let min_68400_45640 = minimum(v(n_68400_45640))
let min_68400_48440 = minimum(v(n_68400_48440))
let min_68400_51240 = minimum(v(n_68400_51240))
let min_68400_54040 = minimum(v(n_68400_54040))
let min_68400_56840 = minimum(v(n_68400_56840))
let min_68400_59640 = minimum(v(n_68400_59640))
let min_68400_62440 = minimum(v(n_68400_62440))
let min_68400_65240 = minimum(v(n_68400_65240))
let min_68400_68040 = minimum(v(n_68400_68040))
let min_68400_70840 = minimum(v(n_68400_70840))
let min_68400_73640 = minimum(v(n_68400_73640))
let min_68400_76440 = minimum(v(n_68400_76440))
let min_68400_79240 = minimum(v(n_68400_79240))
let min_68400_82040 = minimum(v(n_68400_82040))
let min_68400_84840 = minimum(v(n_68400_84840))
let min_68400_87640 = minimum(v(n_68400_87640))
let min_68780_40040 = minimum(v(n_68780_40040))
let min_68780_42840 = minimum(v(n_68780_42840))
let min_68780_45640 = minimum(v(n_68780_45640))
let min_68780_48440 = minimum(v(n_68780_48440))
let min_68780_51240 = minimum(v(n_68780_51240))
let min_68780_54040 = minimum(v(n_68780_54040))
let min_68780_56840 = minimum(v(n_68780_56840))
let min_68780_59640 = minimum(v(n_68780_59640))
let min_68780_62440 = minimum(v(n_68780_62440))
let min_68780_65240 = minimum(v(n_68780_65240))
let min_68780_68040 = minimum(v(n_68780_68040))
let min_68780_70840 = minimum(v(n_68780_70840))
let min_68780_73640 = minimum(v(n_68780_73640))
let min_68780_76440 = minimum(v(n_68780_76440))
let min_68780_79240 = minimum(v(n_68780_79240))
let min_68780_82040 = minimum(v(n_68780_82040))
let min_68780_84840 = minimum(v(n_68780_84840))
let min_68780_87640 = minimum(v(n_68780_87640))
let min_69160_40040 = minimum(v(n_69160_40040))
let min_69160_42840 = minimum(v(n_69160_42840))
let min_69160_45640 = minimum(v(n_69160_45640))
let min_69160_48440 = minimum(v(n_69160_48440))
let min_69160_51240 = minimum(v(n_69160_51240))
let min_69160_54040 = minimum(v(n_69160_54040))
let min_69160_56840 = minimum(v(n_69160_56840))
let min_69160_59640 = minimum(v(n_69160_59640))
let min_69160_62440 = minimum(v(n_69160_62440))
let min_69160_65240 = minimum(v(n_69160_65240))
let min_69160_68040 = minimum(v(n_69160_68040))
let min_69160_70840 = minimum(v(n_69160_70840))
let min_69160_73640 = minimum(v(n_69160_73640))
let min_69160_76440 = minimum(v(n_69160_76440))
let min_69160_79240 = minimum(v(n_69160_79240))
let min_69160_82040 = minimum(v(n_69160_82040))
let min_69160_84840 = minimum(v(n_69160_84840))
let min_69160_87640 = minimum(v(n_69160_87640))
let min_69920_40040 = minimum(v(n_69920_40040))
let min_69920_42840 = minimum(v(n_69920_42840))
let min_69920_45640 = minimum(v(n_69920_45640))
let min_69920_48440 = minimum(v(n_69920_48440))
let min_69920_51240 = minimum(v(n_69920_51240))
let min_69920_54040 = minimum(v(n_69920_54040))
let min_69920_56840 = minimum(v(n_69920_56840))
let min_69920_59640 = minimum(v(n_69920_59640))
let min_69920_62440 = minimum(v(n_69920_62440))
let min_69920_65240 = minimum(v(n_69920_65240))
let min_69920_68040 = minimum(v(n_69920_68040))
let min_69920_70840 = minimum(v(n_69920_70840))
let min_69920_73640 = minimum(v(n_69920_73640))
let min_69920_76440 = minimum(v(n_69920_76440))
let min_69920_79240 = minimum(v(n_69920_79240))
let min_69920_82040 = minimum(v(n_69920_82040))
let min_69920_84840 = minimum(v(n_69920_84840))
let min_69920_87640 = minimum(v(n_69920_87640))
let min_70300_40040 = minimum(v(n_70300_40040))
let min_70300_42840 = minimum(v(n_70300_42840))
let min_70300_45640 = minimum(v(n_70300_45640))
let min_70300_48440 = minimum(v(n_70300_48440))
let min_70300_51240 = minimum(v(n_70300_51240))
let min_70300_54040 = minimum(v(n_70300_54040))
let min_70300_56840 = minimum(v(n_70300_56840))
let min_70300_59640 = minimum(v(n_70300_59640))
let min_70300_62440 = minimum(v(n_70300_62440))
let min_70300_65240 = minimum(v(n_70300_65240))
let min_70300_68040 = minimum(v(n_70300_68040))
let min_70300_70840 = minimum(v(n_70300_70840))
let min_70300_73640 = minimum(v(n_70300_73640))
let min_70300_76440 = minimum(v(n_70300_76440))
let min_70300_79240 = minimum(v(n_70300_79240))
let min_70300_82040 = minimum(v(n_70300_82040))
let min_70300_84840 = minimum(v(n_70300_84840))
let min_70300_87640 = minimum(v(n_70300_87640))
let min_71060_40040 = minimum(v(n_71060_40040))
let min_71060_42840 = minimum(v(n_71060_42840))
let min_71060_45640 = minimum(v(n_71060_45640))
let min_71060_48440 = minimum(v(n_71060_48440))
let min_71060_51240 = minimum(v(n_71060_51240))
let min_71060_54040 = minimum(v(n_71060_54040))
let min_71060_56840 = minimum(v(n_71060_56840))
let min_71060_59640 = minimum(v(n_71060_59640))
let min_71060_62440 = minimum(v(n_71060_62440))
let min_71060_65240 = minimum(v(n_71060_65240))
let min_71060_68040 = minimum(v(n_71060_68040))
let min_71060_70840 = minimum(v(n_71060_70840))
let min_71060_73640 = minimum(v(n_71060_73640))
let min_71060_76440 = minimum(v(n_71060_76440))
let min_71060_79240 = minimum(v(n_71060_79240))
let min_71060_82040 = minimum(v(n_71060_82040))
let min_71060_84840 = minimum(v(n_71060_84840))
let min_71060_87640 = minimum(v(n_71060_87640))
let min_71820_40040 = minimum(v(n_71820_40040))
let min_71820_42840 = minimum(v(n_71820_42840))
let min_71820_45640 = minimum(v(n_71820_45640))
let min_71820_48440 = minimum(v(n_71820_48440))
let min_71820_51240 = minimum(v(n_71820_51240))
let min_71820_54040 = minimum(v(n_71820_54040))
let min_71820_56840 = minimum(v(n_71820_56840))
let min_71820_59640 = minimum(v(n_71820_59640))
let min_71820_62440 = minimum(v(n_71820_62440))
let min_71820_65240 = minimum(v(n_71820_65240))
let min_71820_68040 = minimum(v(n_71820_68040))
let min_71820_70840 = minimum(v(n_71820_70840))
let min_71820_73640 = minimum(v(n_71820_73640))
let min_71820_76440 = minimum(v(n_71820_76440))
let min_71820_79240 = minimum(v(n_71820_79240))
let min_71820_82040 = minimum(v(n_71820_82040))
let min_71820_84840 = minimum(v(n_71820_84840))
let min_71820_87640 = minimum(v(n_71820_87640))
let min_72200_40040 = minimum(v(n_72200_40040))
let min_72200_42840 = minimum(v(n_72200_42840))
let min_72200_45640 = minimum(v(n_72200_45640))
let min_72200_48440 = minimum(v(n_72200_48440))
let min_72200_51240 = minimum(v(n_72200_51240))
let min_72200_54040 = minimum(v(n_72200_54040))
let min_72200_56840 = minimum(v(n_72200_56840))
let min_72200_59640 = minimum(v(n_72200_59640))
let min_72200_62440 = minimum(v(n_72200_62440))
let min_72200_65240 = minimum(v(n_72200_65240))
let min_72200_68040 = minimum(v(n_72200_68040))
let min_72200_70840 = minimum(v(n_72200_70840))
let min_72200_73640 = minimum(v(n_72200_73640))
let min_72200_76440 = minimum(v(n_72200_76440))
let min_72200_79240 = minimum(v(n_72200_79240))
let min_72200_82040 = minimum(v(n_72200_82040))
let min_72200_84840 = minimum(v(n_72200_84840))
let min_72200_87640 = minimum(v(n_72200_87640))
let min_72960_40040 = minimum(v(n_72960_40040))
let min_72960_42840 = minimum(v(n_72960_42840))
let min_72960_45640 = minimum(v(n_72960_45640))
let min_72960_48440 = minimum(v(n_72960_48440))
let min_72960_51240 = minimum(v(n_72960_51240))
let min_72960_54040 = minimum(v(n_72960_54040))
let min_72960_56840 = minimum(v(n_72960_56840))
let min_72960_59640 = minimum(v(n_72960_59640))
let min_72960_62440 = minimum(v(n_72960_62440))
let min_72960_65240 = minimum(v(n_72960_65240))
let min_72960_68040 = minimum(v(n_72960_68040))
let min_72960_70840 = minimum(v(n_72960_70840))
let min_72960_73640 = minimum(v(n_72960_73640))
let min_72960_76440 = minimum(v(n_72960_76440))
let min_72960_79240 = minimum(v(n_72960_79240))
let min_72960_82040 = minimum(v(n_72960_82040))
let min_72960_84840 = minimum(v(n_72960_84840))
let min_72960_87640 = minimum(v(n_72960_87640))
let min_73340_40040 = minimum(v(n_73340_40040))
let min_73340_42840 = minimum(v(n_73340_42840))
let min_73340_45640 = minimum(v(n_73340_45640))
let min_73340_48440 = minimum(v(n_73340_48440))
let min_73340_51240 = minimum(v(n_73340_51240))
let min_73340_54040 = minimum(v(n_73340_54040))
let min_73340_56840 = minimum(v(n_73340_56840))
let min_73340_59640 = minimum(v(n_73340_59640))
let min_73340_62440 = minimum(v(n_73340_62440))
let min_73340_65240 = minimum(v(n_73340_65240))
let min_73340_68040 = minimum(v(n_73340_68040))
let min_73340_70840 = minimum(v(n_73340_70840))
let min_73340_73640 = minimum(v(n_73340_73640))
let min_73340_76440 = minimum(v(n_73340_76440))
let min_73340_79240 = minimum(v(n_73340_79240))
let min_73340_82040 = minimum(v(n_73340_82040))
let min_73340_84840 = minimum(v(n_73340_84840))
let min_73340_87640 = minimum(v(n_73340_87640))
let min_73720_40040 = minimum(v(n_73720_40040))
let min_73720_42840 = minimum(v(n_73720_42840))
let min_73720_45640 = minimum(v(n_73720_45640))
let min_73720_48440 = minimum(v(n_73720_48440))
let min_73720_51240 = minimum(v(n_73720_51240))
let min_73720_54040 = minimum(v(n_73720_54040))
let min_73720_56840 = minimum(v(n_73720_56840))
let min_73720_59640 = minimum(v(n_73720_59640))
let min_73720_62440 = minimum(v(n_73720_62440))
let min_73720_65240 = minimum(v(n_73720_65240))
let min_73720_68040 = minimum(v(n_73720_68040))
let min_73720_70840 = minimum(v(n_73720_70840))
let min_73720_73640 = minimum(v(n_73720_73640))
let min_73720_76440 = minimum(v(n_73720_76440))
let min_73720_79240 = minimum(v(n_73720_79240))
let min_73720_82040 = minimum(v(n_73720_82040))
let min_73720_84840 = minimum(v(n_73720_84840))
let min_73720_87640 = minimum(v(n_73720_87640))
let min_74100_40040 = minimum(v(n_74100_40040))
let min_74100_42840 = minimum(v(n_74100_42840))
let min_74100_45640 = minimum(v(n_74100_45640))
let min_74100_48440 = minimum(v(n_74100_48440))
let min_74100_51240 = minimum(v(n_74100_51240))
let min_74100_54040 = minimum(v(n_74100_54040))
let min_74100_56840 = minimum(v(n_74100_56840))
let min_74100_59640 = minimum(v(n_74100_59640))
let min_74100_62440 = minimum(v(n_74100_62440))
let min_74100_65240 = minimum(v(n_74100_65240))
let min_74100_68040 = minimum(v(n_74100_68040))
let min_74100_70840 = minimum(v(n_74100_70840))
let min_74100_73640 = minimum(v(n_74100_73640))
let min_74100_76440 = minimum(v(n_74100_76440))
let min_74100_79240 = minimum(v(n_74100_79240))
let min_74100_82040 = minimum(v(n_74100_82040))
let min_74100_84840 = minimum(v(n_74100_84840))
let min_74100_87640 = minimum(v(n_74100_87640))
let min_74860_40040 = minimum(v(n_74860_40040))
let min_74860_42840 = minimum(v(n_74860_42840))
let min_74860_45640 = minimum(v(n_74860_45640))
let min_74860_48440 = minimum(v(n_74860_48440))
let min_74860_51240 = minimum(v(n_74860_51240))
let min_74860_54040 = minimum(v(n_74860_54040))
let min_74860_56840 = minimum(v(n_74860_56840))
let min_74860_59640 = minimum(v(n_74860_59640))
let min_74860_62440 = minimum(v(n_74860_62440))
let min_74860_65240 = minimum(v(n_74860_65240))
let min_74860_68040 = minimum(v(n_74860_68040))
let min_74860_70840 = minimum(v(n_74860_70840))
let min_74860_73640 = minimum(v(n_74860_73640))
let min_74860_76440 = minimum(v(n_74860_76440))
let min_74860_79240 = minimum(v(n_74860_79240))
let min_74860_82040 = minimum(v(n_74860_82040))
let min_74860_84840 = minimum(v(n_74860_84840))
let min_74860_87640 = minimum(v(n_74860_87640))
let min_75240_40040 = minimum(v(n_75240_40040))
let min_75240_42840 = minimum(v(n_75240_42840))
let min_75240_45640 = minimum(v(n_75240_45640))
let min_75240_48440 = minimum(v(n_75240_48440))
let min_75240_51240 = minimum(v(n_75240_51240))
let min_75240_54040 = minimum(v(n_75240_54040))
let min_75240_56840 = minimum(v(n_75240_56840))
let min_75240_59640 = minimum(v(n_75240_59640))
let min_75240_62440 = minimum(v(n_75240_62440))
let min_75240_65240 = minimum(v(n_75240_65240))
let min_75240_68040 = minimum(v(n_75240_68040))
let min_75240_70840 = minimum(v(n_75240_70840))
let min_75240_73640 = minimum(v(n_75240_73640))
let min_75240_76440 = minimum(v(n_75240_76440))
let min_75240_79240 = minimum(v(n_75240_79240))
let min_75240_82040 = minimum(v(n_75240_82040))
let min_75240_84840 = minimum(v(n_75240_84840))
let min_75240_87640 = minimum(v(n_75240_87640))
let min_76000_40040 = minimum(v(n_76000_40040))
let min_76000_42840 = minimum(v(n_76000_42840))
let min_76000_45640 = minimum(v(n_76000_45640))
let min_76000_48440 = minimum(v(n_76000_48440))
let min_76000_51240 = minimum(v(n_76000_51240))
let min_76000_54040 = minimum(v(n_76000_54040))
let min_76000_56840 = minimum(v(n_76000_56840))
let min_76000_59640 = minimum(v(n_76000_59640))
let min_76000_62440 = minimum(v(n_76000_62440))
let min_76000_65240 = minimum(v(n_76000_65240))
let min_76000_68040 = minimum(v(n_76000_68040))
let min_76000_70840 = minimum(v(n_76000_70840))
let min_76000_73640 = minimum(v(n_76000_73640))
let min_76000_76440 = minimum(v(n_76000_76440))
let min_76000_79240 = minimum(v(n_76000_79240))
let min_76000_82040 = minimum(v(n_76000_82040))
let min_76000_84840 = minimum(v(n_76000_84840))
let min_76000_87640 = minimum(v(n_76000_87640))
let min_76380_40040 = minimum(v(n_76380_40040))
let min_76380_42840 = minimum(v(n_76380_42840))
let min_76380_45640 = minimum(v(n_76380_45640))
let min_76380_48440 = minimum(v(n_76380_48440))
let min_76380_51240 = minimum(v(n_76380_51240))
let min_76380_54040 = minimum(v(n_76380_54040))
let min_76380_56840 = minimum(v(n_76380_56840))
let min_76380_59640 = minimum(v(n_76380_59640))
let min_76380_62440 = minimum(v(n_76380_62440))
let min_76380_65240 = minimum(v(n_76380_65240))
let min_76380_68040 = minimum(v(n_76380_68040))
let min_76380_70840 = minimum(v(n_76380_70840))
let min_76380_73640 = minimum(v(n_76380_73640))
let min_76380_76440 = minimum(v(n_76380_76440))
let min_76380_79240 = minimum(v(n_76380_79240))
let min_76380_82040 = minimum(v(n_76380_82040))
let min_76380_84840 = minimum(v(n_76380_84840))
let min_76380_87640 = minimum(v(n_76380_87640))
let min_76760_40040 = minimum(v(n_76760_40040))
let min_76760_42840 = minimum(v(n_76760_42840))
let min_76760_45640 = minimum(v(n_76760_45640))
let min_76760_48440 = minimum(v(n_76760_48440))
let min_76760_51240 = minimum(v(n_76760_51240))
let min_76760_54040 = minimum(v(n_76760_54040))
let min_76760_56840 = minimum(v(n_76760_56840))
let min_76760_59640 = minimum(v(n_76760_59640))
let min_76760_62440 = minimum(v(n_76760_62440))
let min_76760_65240 = minimum(v(n_76760_65240))
let min_76760_68040 = minimum(v(n_76760_68040))
let min_76760_70840 = minimum(v(n_76760_70840))
let min_76760_73640 = minimum(v(n_76760_73640))
let min_76760_76440 = minimum(v(n_76760_76440))
let min_76760_79240 = minimum(v(n_76760_79240))
let min_76760_82040 = minimum(v(n_76760_82040))
let min_76760_84840 = minimum(v(n_76760_84840))
let min_76760_87640 = minimum(v(n_76760_87640))
let min_77140_40040 = minimum(v(n_77140_40040))
let min_77140_42840 = minimum(v(n_77140_42840))
let min_77140_45640 = minimum(v(n_77140_45640))
let min_77140_48440 = minimum(v(n_77140_48440))
let min_77140_51240 = minimum(v(n_77140_51240))
let min_77140_54040 = minimum(v(n_77140_54040))
let min_77140_56840 = minimum(v(n_77140_56840))
let min_77140_59640 = minimum(v(n_77140_59640))
let min_77140_62440 = minimum(v(n_77140_62440))
let min_77140_65240 = minimum(v(n_77140_65240))
let min_77140_68040 = minimum(v(n_77140_68040))
let min_77140_70840 = minimum(v(n_77140_70840))
let min_77140_73640 = minimum(v(n_77140_73640))
let min_77140_76440 = minimum(v(n_77140_76440))
let min_77140_79240 = minimum(v(n_77140_79240))
let min_77140_82040 = minimum(v(n_77140_82040))
let min_77140_84840 = minimum(v(n_77140_84840))
let min_77140_87640 = minimum(v(n_77140_87640))
let min_77520_40040 = minimum(v(n_77520_40040))
let min_77520_42840 = minimum(v(n_77520_42840))
let min_77520_45640 = minimum(v(n_77520_45640))
let min_77520_48440 = minimum(v(n_77520_48440))
let min_77520_51240 = minimum(v(n_77520_51240))
let min_77520_54040 = minimum(v(n_77520_54040))
let min_77520_56840 = minimum(v(n_77520_56840))
let min_77520_59640 = minimum(v(n_77520_59640))
let min_77520_62440 = minimum(v(n_77520_62440))
let min_77520_65240 = minimum(v(n_77520_65240))
let min_77520_68040 = minimum(v(n_77520_68040))
let min_77520_70840 = minimum(v(n_77520_70840))
let min_77520_73640 = minimum(v(n_77520_73640))
let min_77520_76440 = minimum(v(n_77520_76440))
let min_77520_79240 = minimum(v(n_77520_79240))
let min_77520_82040 = minimum(v(n_77520_82040))
let min_77520_84840 = minimum(v(n_77520_84840))
let min_77520_87640 = minimum(v(n_77520_87640))
let min_77900_40040 = minimum(v(n_77900_40040))
let min_77900_42840 = minimum(v(n_77900_42840))
let min_77900_45640 = minimum(v(n_77900_45640))
let min_77900_48440 = minimum(v(n_77900_48440))
let min_77900_51240 = minimum(v(n_77900_51240))
let min_77900_54040 = minimum(v(n_77900_54040))
let min_77900_56840 = minimum(v(n_77900_56840))
let min_77900_59640 = minimum(v(n_77900_59640))
let min_77900_62440 = minimum(v(n_77900_62440))
let min_77900_65240 = minimum(v(n_77900_65240))
let min_77900_68040 = minimum(v(n_77900_68040))
let min_77900_70840 = minimum(v(n_77900_70840))
let min_77900_73640 = minimum(v(n_77900_73640))
let min_77900_76440 = minimum(v(n_77900_76440))
let min_77900_79240 = minimum(v(n_77900_79240))
let min_77900_82040 = minimum(v(n_77900_82040))
let min_77900_84840 = minimum(v(n_77900_84840))
let min_77900_87640 = minimum(v(n_77900_87640))
let min_78280_40040 = minimum(v(n_78280_40040))
let min_78280_42840 = minimum(v(n_78280_42840))
let min_78280_45640 = minimum(v(n_78280_45640))
let min_78280_48440 = minimum(v(n_78280_48440))
let min_78280_51240 = minimum(v(n_78280_51240))
let min_78280_54040 = minimum(v(n_78280_54040))
let min_78280_56840 = minimum(v(n_78280_56840))
let min_78280_59640 = minimum(v(n_78280_59640))
let min_78280_62440 = minimum(v(n_78280_62440))
let min_78280_65240 = minimum(v(n_78280_65240))
let min_78280_68040 = minimum(v(n_78280_68040))
let min_78280_70840 = minimum(v(n_78280_70840))
let min_78280_73640 = minimum(v(n_78280_73640))
let min_78280_76440 = minimum(v(n_78280_76440))
let min_78280_79240 = minimum(v(n_78280_79240))
let min_78280_82040 = minimum(v(n_78280_82040))
let min_78280_84840 = minimum(v(n_78280_84840))
let min_78280_87640 = minimum(v(n_78280_87640))
let min_78660_40040 = minimum(v(n_78660_40040))
let min_78660_42840 = minimum(v(n_78660_42840))
let min_78660_45640 = minimum(v(n_78660_45640))
let min_78660_48440 = minimum(v(n_78660_48440))
let min_78660_51240 = minimum(v(n_78660_51240))
let min_78660_54040 = minimum(v(n_78660_54040))
let min_78660_56840 = minimum(v(n_78660_56840))
let min_78660_59640 = minimum(v(n_78660_59640))
let min_78660_62440 = minimum(v(n_78660_62440))
let min_78660_65240 = minimum(v(n_78660_65240))
let min_78660_68040 = minimum(v(n_78660_68040))
let min_78660_70840 = minimum(v(n_78660_70840))
let min_78660_73640 = minimum(v(n_78660_73640))
let min_78660_76440 = minimum(v(n_78660_76440))
let min_78660_79240 = minimum(v(n_78660_79240))
let min_78660_82040 = minimum(v(n_78660_82040))
let min_78660_84840 = minimum(v(n_78660_84840))
let min_78660_87640 = minimum(v(n_78660_87640))
let min_79040_40040 = minimum(v(n_79040_40040))
let min_79040_42840 = minimum(v(n_79040_42840))
let min_79040_45640 = minimum(v(n_79040_45640))
let min_79040_48440 = minimum(v(n_79040_48440))
let min_79040_51240 = minimum(v(n_79040_51240))
let min_79040_54040 = minimum(v(n_79040_54040))
let min_79040_56840 = minimum(v(n_79040_56840))
let min_79040_59640 = minimum(v(n_79040_59640))
let min_79040_62440 = minimum(v(n_79040_62440))
let min_79040_65240 = minimum(v(n_79040_65240))
let min_79040_68040 = minimum(v(n_79040_68040))
let min_79040_70840 = minimum(v(n_79040_70840))
let min_79040_73640 = minimum(v(n_79040_73640))
let min_79040_76440 = minimum(v(n_79040_76440))
let min_79040_79240 = minimum(v(n_79040_79240))
let min_79040_82040 = minimum(v(n_79040_82040))
let min_79040_84840 = minimum(v(n_79040_84840))
let min_79040_87640 = minimum(v(n_79040_87640))
let min_80180_40040 = minimum(v(n_80180_40040))
let min_80180_42840 = minimum(v(n_80180_42840))
let min_80180_45640 = minimum(v(n_80180_45640))
let min_80180_48440 = minimum(v(n_80180_48440))
let min_80180_51240 = minimum(v(n_80180_51240))
let min_80180_54040 = minimum(v(n_80180_54040))
let min_80180_56840 = minimum(v(n_80180_56840))
let min_80180_59640 = minimum(v(n_80180_59640))
let min_80180_62440 = minimum(v(n_80180_62440))
let min_80180_65240 = minimum(v(n_80180_65240))
let min_80180_68040 = minimum(v(n_80180_68040))
let min_80180_70840 = minimum(v(n_80180_70840))
let min_80180_73640 = minimum(v(n_80180_73640))
let min_80180_76440 = minimum(v(n_80180_76440))
let min_80180_79240 = minimum(v(n_80180_79240))
let min_80180_82040 = minimum(v(n_80180_82040))
let min_80180_84840 = minimum(v(n_80180_84840))
let min_80180_87640 = minimum(v(n_80180_87640))
let min_80560_40040 = minimum(v(n_80560_40040))
let min_80560_42840 = minimum(v(n_80560_42840))
let min_80560_45640 = minimum(v(n_80560_45640))
let min_80560_48440 = minimum(v(n_80560_48440))
let min_80560_51240 = minimum(v(n_80560_51240))
let min_80560_54040 = minimum(v(n_80560_54040))
let min_80560_56840 = minimum(v(n_80560_56840))
let min_80560_59640 = minimum(v(n_80560_59640))
let min_80560_62440 = minimum(v(n_80560_62440))
let min_80560_65240 = minimum(v(n_80560_65240))
let min_80560_68040 = minimum(v(n_80560_68040))
let min_80560_70840 = minimum(v(n_80560_70840))
let min_80560_73640 = minimum(v(n_80560_73640))
let min_80560_76440 = minimum(v(n_80560_76440))
let min_80560_79240 = minimum(v(n_80560_79240))
let min_80560_82040 = minimum(v(n_80560_82040))
let min_80560_84840 = minimum(v(n_80560_84840))
let min_80560_87640 = minimum(v(n_80560_87640))
let min_80940_40040 = minimum(v(n_80940_40040))
let min_80940_42840 = minimum(v(n_80940_42840))
let min_80940_45640 = minimum(v(n_80940_45640))
let min_80940_48440 = minimum(v(n_80940_48440))
let min_80940_51240 = minimum(v(n_80940_51240))
let min_80940_54040 = minimum(v(n_80940_54040))
let min_80940_56840 = minimum(v(n_80940_56840))
let min_80940_59640 = minimum(v(n_80940_59640))
let min_80940_62440 = minimum(v(n_80940_62440))
let min_80940_65240 = minimum(v(n_80940_65240))
let min_80940_68040 = minimum(v(n_80940_68040))
let min_80940_70840 = minimum(v(n_80940_70840))
let min_80940_73640 = minimum(v(n_80940_73640))
let min_80940_76440 = minimum(v(n_80940_76440))
let min_80940_79240 = minimum(v(n_80940_79240))
let min_80940_82040 = minimum(v(n_80940_82040))
let min_80940_84840 = minimum(v(n_80940_84840))
let min_80940_87640 = minimum(v(n_80940_87640))
let min_81700_40040 = minimum(v(n_81700_40040))
let min_81700_42840 = minimum(v(n_81700_42840))
let min_81700_45640 = minimum(v(n_81700_45640))
let min_81700_48440 = minimum(v(n_81700_48440))
let min_81700_51240 = minimum(v(n_81700_51240))
let min_81700_54040 = minimum(v(n_81700_54040))
let min_81700_56840 = minimum(v(n_81700_56840))
let min_81700_59640 = minimum(v(n_81700_59640))
let min_81700_62440 = minimum(v(n_81700_62440))
let min_81700_65240 = minimum(v(n_81700_65240))
let min_81700_68040 = minimum(v(n_81700_68040))
let min_81700_70840 = minimum(v(n_81700_70840))
let min_81700_73640 = minimum(v(n_81700_73640))
let min_81700_76440 = minimum(v(n_81700_76440))
let min_81700_79240 = minimum(v(n_81700_79240))
let min_81700_82040 = minimum(v(n_81700_82040))
let min_81700_84840 = minimum(v(n_81700_84840))
let min_81700_87640 = minimum(v(n_81700_87640))
let min_82080_40040 = minimum(v(n_82080_40040))
let min_82080_42840 = minimum(v(n_82080_42840))
let min_82080_45640 = minimum(v(n_82080_45640))
let min_82080_48440 = minimum(v(n_82080_48440))
let min_82080_51240 = minimum(v(n_82080_51240))
let min_82080_54040 = minimum(v(n_82080_54040))
let min_82080_56840 = minimum(v(n_82080_56840))
let min_82080_59640 = minimum(v(n_82080_59640))
let min_82080_62440 = minimum(v(n_82080_62440))
let min_82080_65240 = minimum(v(n_82080_65240))
let min_82080_68040 = minimum(v(n_82080_68040))
let min_82080_70840 = minimum(v(n_82080_70840))
let min_82080_73640 = minimum(v(n_82080_73640))
let min_82080_76440 = minimum(v(n_82080_76440))
let min_82080_79240 = minimum(v(n_82080_79240))
let min_82080_82040 = minimum(v(n_82080_82040))
let min_82080_84840 = minimum(v(n_82080_84840))
let min_82080_87640 = minimum(v(n_82080_87640))
let min_83220_40040 = minimum(v(n_83220_40040))
let min_83220_42840 = minimum(v(n_83220_42840))
let min_83220_45640 = minimum(v(n_83220_45640))
let min_83220_48440 = minimum(v(n_83220_48440))
let min_83220_51240 = minimum(v(n_83220_51240))
let min_83220_54040 = minimum(v(n_83220_54040))
let min_83220_56840 = minimum(v(n_83220_56840))
let min_83220_59640 = minimum(v(n_83220_59640))
let min_83220_62440 = minimum(v(n_83220_62440))
let min_83220_65240 = minimum(v(n_83220_65240))
let min_83220_68040 = minimum(v(n_83220_68040))
let min_83220_70840 = minimum(v(n_83220_70840))
let min_83220_73640 = minimum(v(n_83220_73640))
let min_83220_76440 = minimum(v(n_83220_76440))
let min_83220_79240 = minimum(v(n_83220_79240))
let min_83220_82040 = minimum(v(n_83220_82040))
let min_83220_84840 = minimum(v(n_83220_84840))
let min_83220_87640 = minimum(v(n_83220_87640))
let min_83600_40040 = minimum(v(n_83600_40040))
let min_83600_42840 = minimum(v(n_83600_42840))
let min_83600_45640 = minimum(v(n_83600_45640))
let min_83600_48440 = minimum(v(n_83600_48440))
let min_83600_51240 = minimum(v(n_83600_51240))
let min_83600_54040 = minimum(v(n_83600_54040))
let min_83600_56840 = minimum(v(n_83600_56840))
let min_83600_59640 = minimum(v(n_83600_59640))
let min_83600_62440 = minimum(v(n_83600_62440))
let min_83600_65240 = minimum(v(n_83600_65240))
let min_83600_68040 = minimum(v(n_83600_68040))
let min_83600_70840 = minimum(v(n_83600_70840))
let min_83600_73640 = minimum(v(n_83600_73640))
let min_83600_76440 = minimum(v(n_83600_76440))
let min_83600_79240 = minimum(v(n_83600_79240))
let min_83600_82040 = minimum(v(n_83600_82040))
let min_83600_84840 = minimum(v(n_83600_84840))
let min_83600_87640 = minimum(v(n_83600_87640))
let min_84740_40040 = minimum(v(n_84740_40040))
let min_84740_42840 = minimum(v(n_84740_42840))
let min_84740_45640 = minimum(v(n_84740_45640))
let min_84740_48440 = minimum(v(n_84740_48440))
let min_84740_51240 = minimum(v(n_84740_51240))
let min_84740_54040 = minimum(v(n_84740_54040))
let min_84740_56840 = minimum(v(n_84740_56840))
let min_84740_59640 = minimum(v(n_84740_59640))
let min_84740_62440 = minimum(v(n_84740_62440))
let min_84740_65240 = minimum(v(n_84740_65240))
let min_84740_68040 = minimum(v(n_84740_68040))
let min_84740_70840 = minimum(v(n_84740_70840))
let min_84740_73640 = minimum(v(n_84740_73640))
let min_84740_76440 = minimum(v(n_84740_76440))
let min_84740_79240 = minimum(v(n_84740_79240))
let min_84740_82040 = minimum(v(n_84740_82040))
let min_84740_84840 = minimum(v(n_84740_84840))
let min_84740_87640 = minimum(v(n_84740_87640))
let min_85120_40040 = minimum(v(n_85120_40040))
let min_85120_42840 = minimum(v(n_85120_42840))
let min_85120_45640 = minimum(v(n_85120_45640))
let min_85120_48440 = minimum(v(n_85120_48440))
let min_85120_51240 = minimum(v(n_85120_51240))
let min_85120_54040 = minimum(v(n_85120_54040))
let min_85120_56840 = minimum(v(n_85120_56840))
let min_85120_59640 = minimum(v(n_85120_59640))
let min_85120_62440 = minimum(v(n_85120_62440))
let min_85120_65240 = minimum(v(n_85120_65240))
let min_85120_68040 = minimum(v(n_85120_68040))
let min_85120_70840 = minimum(v(n_85120_70840))
let min_85120_73640 = minimum(v(n_85120_73640))
let min_85120_76440 = minimum(v(n_85120_76440))
let min_85120_79240 = minimum(v(n_85120_79240))
let min_85120_82040 = minimum(v(n_85120_82040))
let min_85120_84840 = minimum(v(n_85120_84840))
let min_85120_87640 = minimum(v(n_85120_87640))
let min_85500_40040 = minimum(v(n_85500_40040))
let min_85500_42840 = minimum(v(n_85500_42840))
let min_85500_45640 = minimum(v(n_85500_45640))
let min_85500_48440 = minimum(v(n_85500_48440))
let min_85500_51240 = minimum(v(n_85500_51240))
let min_85500_54040 = minimum(v(n_85500_54040))
let min_85500_56840 = minimum(v(n_85500_56840))
let min_85500_59640 = minimum(v(n_85500_59640))
let min_85500_62440 = minimum(v(n_85500_62440))
let min_85500_65240 = minimum(v(n_85500_65240))
let min_85500_68040 = minimum(v(n_85500_68040))
let min_85500_70840 = minimum(v(n_85500_70840))
let min_85500_73640 = minimum(v(n_85500_73640))
let min_85500_76440 = minimum(v(n_85500_76440))
let min_85500_79240 = minimum(v(n_85500_79240))
let min_85500_82040 = minimum(v(n_85500_82040))
let min_85500_84840 = minimum(v(n_85500_84840))
let min_85500_87640 = minimum(v(n_85500_87640))
let min_85880_40040 = minimum(v(n_85880_40040))
let min_85880_42840 = minimum(v(n_85880_42840))
let min_85880_45640 = minimum(v(n_85880_45640))
let min_85880_48440 = minimum(v(n_85880_48440))
let min_85880_51240 = minimum(v(n_85880_51240))
let min_85880_54040 = minimum(v(n_85880_54040))
let min_85880_56840 = minimum(v(n_85880_56840))
let min_85880_59640 = minimum(v(n_85880_59640))
let min_85880_62440 = minimum(v(n_85880_62440))
let min_85880_65240 = minimum(v(n_85880_65240))
let min_85880_68040 = minimum(v(n_85880_68040))
let min_85880_70840 = minimum(v(n_85880_70840))
let min_85880_73640 = minimum(v(n_85880_73640))
let min_85880_76440 = minimum(v(n_85880_76440))
let min_85880_79240 = minimum(v(n_85880_79240))
let min_85880_82040 = minimum(v(n_85880_82040))
let min_85880_84840 = minimum(v(n_85880_84840))
let min_85880_87640 = minimum(v(n_85880_87640))
let min_86260_40040 = minimum(v(n_86260_40040))
let min_86260_42840 = minimum(v(n_86260_42840))
let min_86260_45640 = minimum(v(n_86260_45640))
let min_86260_48440 = minimum(v(n_86260_48440))
let min_86260_51240 = minimum(v(n_86260_51240))
let min_86260_54040 = minimum(v(n_86260_54040))
let min_86260_56840 = minimum(v(n_86260_56840))
let min_86260_59640 = minimum(v(n_86260_59640))
let min_86260_62440 = minimum(v(n_86260_62440))
let min_86260_65240 = minimum(v(n_86260_65240))
let min_86260_68040 = minimum(v(n_86260_68040))
let min_86260_70840 = minimum(v(n_86260_70840))
let min_86260_73640 = minimum(v(n_86260_73640))
let min_86260_76440 = minimum(v(n_86260_76440))
let min_86260_79240 = minimum(v(n_86260_79240))
let min_86260_82040 = minimum(v(n_86260_82040))
let min_86260_84840 = minimum(v(n_86260_84840))
let min_86260_87640 = minimum(v(n_86260_87640))
let min_87020_40040 = minimum(v(n_87020_40040))
let min_87020_42840 = minimum(v(n_87020_42840))
let min_87020_45640 = minimum(v(n_87020_45640))
let min_87020_48440 = minimum(v(n_87020_48440))
let min_87020_51240 = minimum(v(n_87020_51240))
let min_87020_54040 = minimum(v(n_87020_54040))
let min_87020_56840 = minimum(v(n_87020_56840))
let min_87020_59640 = minimum(v(n_87020_59640))
let min_87020_62440 = minimum(v(n_87020_62440))
let min_87020_65240 = minimum(v(n_87020_65240))
let min_87020_68040 = minimum(v(n_87020_68040))
let min_87020_70840 = minimum(v(n_87020_70840))
let min_87020_73640 = minimum(v(n_87020_73640))
let min_87020_76440 = minimum(v(n_87020_76440))
let min_87020_79240 = minimum(v(n_87020_79240))
let min_87020_82040 = minimum(v(n_87020_82040))
let min_87020_84840 = minimum(v(n_87020_84840))
let min_87020_87640 = minimum(v(n_87020_87640))
let min_87400_40040 = minimum(v(n_87400_40040))
let min_87400_42840 = minimum(v(n_87400_42840))
let min_87400_45640 = minimum(v(n_87400_45640))
let min_87400_48440 = minimum(v(n_87400_48440))
let min_87400_51240 = minimum(v(n_87400_51240))
let min_87400_54040 = minimum(v(n_87400_54040))
let min_87400_56840 = minimum(v(n_87400_56840))
let min_87400_59640 = minimum(v(n_87400_59640))
let min_87400_62440 = minimum(v(n_87400_62440))
let min_87400_65240 = minimum(v(n_87400_65240))
let min_87400_68040 = minimum(v(n_87400_68040))
let min_87400_70840 = minimum(v(n_87400_70840))
let min_87400_73640 = minimum(v(n_87400_73640))
let min_87400_76440 = minimum(v(n_87400_76440))
let min_87400_79240 = minimum(v(n_87400_79240))
let min_87400_82040 = minimum(v(n_87400_82040))
let min_87400_84840 = minimum(v(n_87400_84840))
let min_87400_87640 = minimum(v(n_87400_87640))
let min_87780_40040 = minimum(v(n_87780_40040))
let min_87780_42840 = minimum(v(n_87780_42840))
let min_87780_45640 = minimum(v(n_87780_45640))
let min_87780_48440 = minimum(v(n_87780_48440))
let min_87780_51240 = minimum(v(n_87780_51240))
let min_87780_54040 = minimum(v(n_87780_54040))
let min_87780_56840 = minimum(v(n_87780_56840))
let min_87780_59640 = minimum(v(n_87780_59640))
let min_87780_62440 = minimum(v(n_87780_62440))
let min_87780_65240 = minimum(v(n_87780_65240))
let min_87780_68040 = minimum(v(n_87780_68040))
let min_87780_70840 = minimum(v(n_87780_70840))
let min_87780_73640 = minimum(v(n_87780_73640))
let min_87780_76440 = minimum(v(n_87780_76440))
let min_87780_79240 = minimum(v(n_87780_79240))
let min_87780_82040 = minimum(v(n_87780_82040))
let min_87780_84840 = minimum(v(n_87780_84840))
let min_87780_87640 = minimum(v(n_87780_87640))
let min_88160_40040 = minimum(v(n_88160_40040))
let min_88160_42840 = minimum(v(n_88160_42840))
let min_88160_45640 = minimum(v(n_88160_45640))
let min_88160_48440 = minimum(v(n_88160_48440))
let min_88160_51240 = minimum(v(n_88160_51240))
let min_88160_54040 = minimum(v(n_88160_54040))
let min_88160_56840 = minimum(v(n_88160_56840))
let min_88160_59640 = minimum(v(n_88160_59640))
let min_88160_62440 = minimum(v(n_88160_62440))
let min_88160_65240 = minimum(v(n_88160_65240))
let min_88160_68040 = minimum(v(n_88160_68040))
let min_88160_70840 = minimum(v(n_88160_70840))
let min_88160_73640 = minimum(v(n_88160_73640))
let min_88160_76440 = minimum(v(n_88160_76440))
let min_88160_79240 = minimum(v(n_88160_79240))
let min_88160_82040 = minimum(v(n_88160_82040))
let min_88160_84840 = minimum(v(n_88160_84840))
let min_88160_87640 = minimum(v(n_88160_87640))
let min_88540_40040 = minimum(v(n_88540_40040))
let min_88540_42840 = minimum(v(n_88540_42840))
let min_88540_45640 = minimum(v(n_88540_45640))
let min_88540_48440 = minimum(v(n_88540_48440))
let min_88540_51240 = minimum(v(n_88540_51240))
let min_88540_54040 = minimum(v(n_88540_54040))
let min_88540_56840 = minimum(v(n_88540_56840))
let min_88540_59640 = minimum(v(n_88540_59640))
let min_88540_62440 = minimum(v(n_88540_62440))
let min_88540_65240 = minimum(v(n_88540_65240))
let min_88540_68040 = minimum(v(n_88540_68040))
let min_88540_70840 = minimum(v(n_88540_70840))
let min_88540_73640 = minimum(v(n_88540_73640))
let min_88540_76440 = minimum(v(n_88540_76440))
let min_88540_79240 = minimum(v(n_88540_79240))
let min_88540_82040 = minimum(v(n_88540_82040))
let min_88540_84840 = minimum(v(n_88540_84840))
let min_88540_87640 = minimum(v(n_88540_87640))
let min_88920_40040 = minimum(v(n_88920_40040))
let min_88920_42840 = minimum(v(n_88920_42840))
let min_88920_45640 = minimum(v(n_88920_45640))
let min_88920_48440 = minimum(v(n_88920_48440))
let min_88920_51240 = minimum(v(n_88920_51240))
let min_88920_54040 = minimum(v(n_88920_54040))
let min_88920_56840 = minimum(v(n_88920_56840))
let min_88920_59640 = minimum(v(n_88920_59640))
let min_88920_62440 = minimum(v(n_88920_62440))
let min_88920_65240 = minimum(v(n_88920_65240))
let min_88920_68040 = minimum(v(n_88920_68040))
let min_88920_70840 = minimum(v(n_88920_70840))
let min_88920_73640 = minimum(v(n_88920_73640))
let min_88920_76440 = minimum(v(n_88920_76440))
let min_88920_79240 = minimum(v(n_88920_79240))
let min_88920_82040 = minimum(v(n_88920_82040))
let min_88920_84840 = minimum(v(n_88920_84840))
let min_88920_87640 = minimum(v(n_88920_87640))
let min_89300_40040 = minimum(v(n_89300_40040))
let min_89300_42840 = minimum(v(n_89300_42840))
let min_89300_45640 = minimum(v(n_89300_45640))
let min_89300_48440 = minimum(v(n_89300_48440))
let min_89300_51240 = minimum(v(n_89300_51240))
let min_89300_54040 = minimum(v(n_89300_54040))
let min_89300_56840 = minimum(v(n_89300_56840))
let min_89300_59640 = minimum(v(n_89300_59640))
let min_89300_62440 = minimum(v(n_89300_62440))
let min_89300_65240 = minimum(v(n_89300_65240))
let min_89300_68040 = minimum(v(n_89300_68040))
let min_89300_70840 = minimum(v(n_89300_70840))
let min_89300_73640 = minimum(v(n_89300_73640))
let min_89300_76440 = minimum(v(n_89300_76440))
let min_89300_79240 = minimum(v(n_89300_79240))
let min_89300_82040 = minimum(v(n_89300_82040))
let min_89300_84840 = minimum(v(n_89300_84840))
let min_89300_87640 = minimum(v(n_89300_87640))
let min_90060_40040 = minimum(v(n_90060_40040))
let min_90060_42840 = minimum(v(n_90060_42840))
let min_90060_45640 = minimum(v(n_90060_45640))
let min_90060_48440 = minimum(v(n_90060_48440))
let min_90060_51240 = minimum(v(n_90060_51240))
let min_90060_54040 = minimum(v(n_90060_54040))
let min_90060_56840 = minimum(v(n_90060_56840))
let min_90060_59640 = minimum(v(n_90060_59640))
let min_90060_62440 = minimum(v(n_90060_62440))
let min_90060_65240 = minimum(v(n_90060_65240))
let min_90060_68040 = minimum(v(n_90060_68040))
let min_90060_70840 = minimum(v(n_90060_70840))
let min_90060_73640 = minimum(v(n_90060_73640))
let min_90060_76440 = minimum(v(n_90060_76440))
let min_90060_79240 = minimum(v(n_90060_79240))
let min_90060_82040 = minimum(v(n_90060_82040))
let min_90060_84840 = minimum(v(n_90060_84840))
let min_90060_87640 = minimum(v(n_90060_87640))
let min_90440_40040 = minimum(v(n_90440_40040))
let min_90440_42840 = minimum(v(n_90440_42840))
let min_90440_45640 = minimum(v(n_90440_45640))
let min_90440_48440 = minimum(v(n_90440_48440))
let min_90440_51240 = minimum(v(n_90440_51240))
let min_90440_54040 = minimum(v(n_90440_54040))
let min_90440_56840 = minimum(v(n_90440_56840))
let min_90440_59640 = minimum(v(n_90440_59640))
let min_90440_62440 = minimum(v(n_90440_62440))
let min_90440_65240 = minimum(v(n_90440_65240))
let min_90440_68040 = minimum(v(n_90440_68040))
let min_90440_70840 = minimum(v(n_90440_70840))
let min_90440_73640 = minimum(v(n_90440_73640))
let min_90440_76440 = minimum(v(n_90440_76440))
let min_90440_79240 = minimum(v(n_90440_79240))
let min_90440_82040 = minimum(v(n_90440_82040))
let min_90440_84840 = minimum(v(n_90440_84840))
let min_90440_87640 = minimum(v(n_90440_87640))
let min_90820_40040 = minimum(v(n_90820_40040))
let min_90820_42840 = minimum(v(n_90820_42840))
let min_90820_45640 = minimum(v(n_90820_45640))
let min_90820_48440 = minimum(v(n_90820_48440))
let min_90820_51240 = minimum(v(n_90820_51240))
let min_90820_54040 = minimum(v(n_90820_54040))
let min_90820_56840 = minimum(v(n_90820_56840))
let min_90820_59640 = minimum(v(n_90820_59640))
let min_90820_62440 = minimum(v(n_90820_62440))
let min_90820_65240 = minimum(v(n_90820_65240))
let min_90820_68040 = minimum(v(n_90820_68040))
let min_90820_70840 = minimum(v(n_90820_70840))
let min_90820_73640 = minimum(v(n_90820_73640))
let min_90820_76440 = minimum(v(n_90820_76440))
let min_90820_79240 = minimum(v(n_90820_79240))
let min_90820_82040 = minimum(v(n_90820_82040))
let min_90820_84840 = minimum(v(n_90820_84840))
let min_90820_87640 = minimum(v(n_90820_87640))
let min_91200_40040 = minimum(v(n_91200_40040))
let min_91200_42840 = minimum(v(n_91200_42840))
let min_91200_45640 = minimum(v(n_91200_45640))
let min_91200_48440 = minimum(v(n_91200_48440))
let min_91200_51240 = minimum(v(n_91200_51240))
let min_91200_54040 = minimum(v(n_91200_54040))
let min_91200_56840 = minimum(v(n_91200_56840))
let min_91200_59640 = minimum(v(n_91200_59640))
let min_91200_62440 = minimum(v(n_91200_62440))
let min_91200_65240 = minimum(v(n_91200_65240))
let min_91200_68040 = minimum(v(n_91200_68040))
let min_91200_70840 = minimum(v(n_91200_70840))
let min_91200_73640 = minimum(v(n_91200_73640))
let min_91200_76440 = minimum(v(n_91200_76440))
let min_91200_79240 = minimum(v(n_91200_79240))
let min_91200_82040 = minimum(v(n_91200_82040))
let min_91200_84840 = minimum(v(n_91200_84840))
let min_91200_87640 = minimum(v(n_91200_87640))
let min_91580_40040 = minimum(v(n_91580_40040))
let min_91580_42840 = minimum(v(n_91580_42840))
let min_91580_45640 = minimum(v(n_91580_45640))
let min_91580_48440 = minimum(v(n_91580_48440))
let min_91580_51240 = minimum(v(n_91580_51240))
let min_91580_54040 = minimum(v(n_91580_54040))
let min_91580_56840 = minimum(v(n_91580_56840))
let min_91580_59640 = minimum(v(n_91580_59640))
let min_91580_62440 = minimum(v(n_91580_62440))
let min_91580_65240 = minimum(v(n_91580_65240))
let min_91580_68040 = minimum(v(n_91580_68040))
let min_91580_70840 = minimum(v(n_91580_70840))
let min_91580_73640 = minimum(v(n_91580_73640))
let min_91580_76440 = minimum(v(n_91580_76440))
let min_91580_79240 = minimum(v(n_91580_79240))
let min_91580_82040 = minimum(v(n_91580_82040))
let min_91580_84840 = minimum(v(n_91580_84840))
let min_91580_87640 = minimum(v(n_91580_87640))
let min_91960_40040 = minimum(v(n_91960_40040))
let min_91960_42840 = minimum(v(n_91960_42840))
let min_91960_45640 = minimum(v(n_91960_45640))
let min_91960_48440 = minimum(v(n_91960_48440))
let min_91960_51240 = minimum(v(n_91960_51240))
let min_91960_54040 = minimum(v(n_91960_54040))
let min_91960_56840 = minimum(v(n_91960_56840))
let min_91960_59640 = minimum(v(n_91960_59640))
let min_91960_62440 = minimum(v(n_91960_62440))
let min_91960_65240 = minimum(v(n_91960_65240))
let min_91960_68040 = minimum(v(n_91960_68040))
let min_91960_70840 = minimum(v(n_91960_70840))
let min_91960_73640 = minimum(v(n_91960_73640))
let min_91960_76440 = minimum(v(n_91960_76440))
let min_91960_79240 = minimum(v(n_91960_79240))
let min_91960_82040 = minimum(v(n_91960_82040))
let min_91960_84840 = minimum(v(n_91960_84840))
let min_91960_87640 = minimum(v(n_91960_87640))
let min_92340_40040 = minimum(v(n_92340_40040))
let min_92340_42840 = minimum(v(n_92340_42840))
let min_92340_45640 = minimum(v(n_92340_45640))
let min_92340_48440 = minimum(v(n_92340_48440))
let min_92340_51240 = minimum(v(n_92340_51240))
let min_92340_54040 = minimum(v(n_92340_54040))
let min_92340_56840 = minimum(v(n_92340_56840))
let min_92340_59640 = minimum(v(n_92340_59640))
let min_92340_62440 = minimum(v(n_92340_62440))
let min_92340_65240 = minimum(v(n_92340_65240))
let min_92340_68040 = minimum(v(n_92340_68040))
let min_92340_70840 = minimum(v(n_92340_70840))
let min_92340_73640 = minimum(v(n_92340_73640))
let min_92340_76440 = minimum(v(n_92340_76440))
let min_92340_79240 = minimum(v(n_92340_79240))
let min_92340_82040 = minimum(v(n_92340_82040))
let min_92340_84840 = minimum(v(n_92340_84840))
let min_92340_87640 = minimum(v(n_92340_87640))
let min_92720_40040 = minimum(v(n_92720_40040))
let min_92720_42840 = minimum(v(n_92720_42840))
let min_92720_45640 = minimum(v(n_92720_45640))
let min_92720_48440 = minimum(v(n_92720_48440))
let min_92720_51240 = minimum(v(n_92720_51240))
let min_92720_54040 = minimum(v(n_92720_54040))
let min_92720_56840 = minimum(v(n_92720_56840))
let min_92720_59640 = minimum(v(n_92720_59640))
let min_92720_62440 = minimum(v(n_92720_62440))
let min_92720_65240 = minimum(v(n_92720_65240))
let min_92720_68040 = minimum(v(n_92720_68040))
let min_92720_70840 = minimum(v(n_92720_70840))
let min_92720_73640 = minimum(v(n_92720_73640))
let min_92720_76440 = minimum(v(n_92720_76440))
let min_92720_79240 = minimum(v(n_92720_79240))
let min_92720_82040 = minimum(v(n_92720_82040))
let min_92720_84840 = minimum(v(n_92720_84840))
let min_92720_87640 = minimum(v(n_92720_87640))
let min_93100_40040 = minimum(v(n_93100_40040))
let min_93100_42840 = minimum(v(n_93100_42840))
let min_93100_45640 = minimum(v(n_93100_45640))
let min_93100_48440 = minimum(v(n_93100_48440))
let min_93100_51240 = minimum(v(n_93100_51240))
let min_93100_54040 = minimum(v(n_93100_54040))
let min_93100_56840 = minimum(v(n_93100_56840))
let min_93100_59640 = minimum(v(n_93100_59640))
let min_93100_62440 = minimum(v(n_93100_62440))
let min_93100_65240 = minimum(v(n_93100_65240))
let min_93100_68040 = minimum(v(n_93100_68040))
let min_93100_70840 = minimum(v(n_93100_70840))
let min_93100_73640 = minimum(v(n_93100_73640))
let min_93100_76440 = minimum(v(n_93100_76440))
let min_93100_79240 = minimum(v(n_93100_79240))
let min_93100_82040 = minimum(v(n_93100_82040))
let min_93100_84840 = minimum(v(n_93100_84840))
let min_93100_87640 = minimum(v(n_93100_87640))
let min_93480_40040 = minimum(v(n_93480_40040))
let min_93480_42840 = minimum(v(n_93480_42840))
let min_93480_45640 = minimum(v(n_93480_45640))
let min_93480_48440 = minimum(v(n_93480_48440))
let min_93480_51240 = minimum(v(n_93480_51240))
let min_93480_54040 = minimum(v(n_93480_54040))
let min_93480_56840 = minimum(v(n_93480_56840))
let min_93480_59640 = minimum(v(n_93480_59640))
let min_93480_62440 = minimum(v(n_93480_62440))
let min_93480_65240 = minimum(v(n_93480_65240))
let min_93480_68040 = minimum(v(n_93480_68040))
let min_93480_70840 = minimum(v(n_93480_70840))
let min_93480_73640 = minimum(v(n_93480_73640))
let min_93480_76440 = minimum(v(n_93480_76440))
let min_93480_79240 = minimum(v(n_93480_79240))
let min_93480_82040 = minimum(v(n_93480_82040))
let min_93480_84840 = minimum(v(n_93480_84840))
let min_93480_87640 = minimum(v(n_93480_87640))
* now write(append) all minimums to a file. ">>" means append:
print min_40280_40040 >> minimums
print min_40280_42840 >> minimums
print min_40280_45640 >> minimums
print min_40280_48440 >> minimums
print min_40280_51240 >> minimums
print min_40280_54040 >> minimums
print min_40280_56840 >> minimums
print min_40280_59640 >> minimums
print min_40280_62440 >> minimums
print min_40280_65240 >> minimums
print min_40280_68040 >> minimums
print min_40280_70840 >> minimums
print min_40280_73640 >> minimums
print min_40280_76440 >> minimums
print min_40280_79240 >> minimums
print min_40280_82040 >> minimums
print min_40280_84840 >> minimums
print min_40280_87640 >> minimums
print min_40660_40040 >> minimums
print min_40660_42840 >> minimums
print min_40660_45640 >> minimums
print min_40660_48440 >> minimums
print min_40660_51240 >> minimums
print min_40660_54040 >> minimums
print min_40660_56840 >> minimums
print min_40660_59640 >> minimums
print min_40660_62440 >> minimums
print min_40660_65240 >> minimums
print min_40660_68040 >> minimums
print min_40660_70840 >> minimums
print min_40660_73640 >> minimums
print min_40660_76440 >> minimums
print min_40660_79240 >> minimums
print min_40660_82040 >> minimums
print min_40660_84840 >> minimums
print min_40660_87640 >> minimums
print min_41420_40040 >> minimums
print min_41420_42840 >> minimums
print min_41420_45640 >> minimums
print min_41420_48440 >> minimums
print min_41420_51240 >> minimums
print min_41420_54040 >> minimums
print min_41420_56840 >> minimums
print min_41420_59640 >> minimums
print min_41420_62440 >> minimums
print min_41420_65240 >> minimums
print min_41420_68040 >> minimums
print min_41420_70840 >> minimums
print min_41420_73640 >> minimums
print min_41420_76440 >> minimums
print min_41420_79240 >> minimums
print min_41420_82040 >> minimums
print min_41420_84840 >> minimums
print min_41420_87640 >> minimums
print min_41800_40040 >> minimums
print min_41800_42840 >> minimums
print min_41800_45640 >> minimums
print min_41800_48440 >> minimums
print min_41800_51240 >> minimums
print min_41800_54040 >> minimums
print min_41800_56840 >> minimums
print min_41800_59640 >> minimums
print min_41800_62440 >> minimums
print min_41800_65240 >> minimums
print min_41800_68040 >> minimums
print min_41800_70840 >> minimums
print min_41800_73640 >> minimums
print min_41800_76440 >> minimums
print min_41800_79240 >> minimums
print min_41800_82040 >> minimums
print min_41800_84840 >> minimums
print min_41800_87640 >> minimums
print min_42180_40040 >> minimums
print min_42180_42840 >> minimums
print min_42180_45640 >> minimums
print min_42180_48440 >> minimums
print min_42180_51240 >> minimums
print min_42180_54040 >> minimums
print min_42180_56840 >> minimums
print min_42180_59640 >> minimums
print min_42180_62440 >> minimums
print min_42180_65240 >> minimums
print min_42180_68040 >> minimums
print min_42180_70840 >> minimums
print min_42180_73640 >> minimums
print min_42180_76440 >> minimums
print min_42180_79240 >> minimums
print min_42180_82040 >> minimums
print min_42180_84840 >> minimums
print min_42180_87640 >> minimums
print min_42940_40040 >> minimums
print min_42940_42840 >> minimums
print min_42940_45640 >> minimums
print min_42940_48440 >> minimums
print min_42940_51240 >> minimums
print min_42940_54040 >> minimums
print min_42940_56840 >> minimums
print min_42940_59640 >> minimums
print min_42940_62440 >> minimums
print min_42940_65240 >> minimums
print min_42940_68040 >> minimums
print min_42940_70840 >> minimums
print min_42940_73640 >> minimums
print min_42940_76440 >> minimums
print min_42940_79240 >> minimums
print min_42940_82040 >> minimums
print min_42940_84840 >> minimums
print min_42940_87640 >> minimums
print min_43320_40040 >> minimums
print min_43320_42840 >> minimums
print min_43320_45640 >> minimums
print min_43320_48440 >> minimums
print min_43320_51240 >> minimums
print min_43320_54040 >> minimums
print min_43320_56840 >> minimums
print min_43320_59640 >> minimums
print min_43320_62440 >> minimums
print min_43320_65240 >> minimums
print min_43320_68040 >> minimums
print min_43320_70840 >> minimums
print min_43320_73640 >> minimums
print min_43320_76440 >> minimums
print min_43320_79240 >> minimums
print min_43320_82040 >> minimums
print min_43320_84840 >> minimums
print min_43320_87640 >> minimums
print min_43700_40040 >> minimums
print min_43700_42840 >> minimums
print min_43700_45640 >> minimums
print min_43700_48440 >> minimums
print min_43700_51240 >> minimums
print min_43700_54040 >> minimums
print min_43700_56840 >> minimums
print min_43700_59640 >> minimums
print min_43700_62440 >> minimums
print min_43700_65240 >> minimums
print min_43700_68040 >> minimums
print min_43700_70840 >> minimums
print min_43700_73640 >> minimums
print min_43700_76440 >> minimums
print min_43700_79240 >> minimums
print min_43700_82040 >> minimums
print min_43700_84840 >> minimums
print min_43700_87640 >> minimums
print min_44080_40040 >> minimums
print min_44080_42840 >> minimums
print min_44080_45640 >> minimums
print min_44080_48440 >> minimums
print min_44080_51240 >> minimums
print min_44080_54040 >> minimums
print min_44080_56840 >> minimums
print min_44080_59640 >> minimums
print min_44080_62440 >> minimums
print min_44080_65240 >> minimums
print min_44080_68040 >> minimums
print min_44080_70840 >> minimums
print min_44080_73640 >> minimums
print min_44080_76440 >> minimums
print min_44080_79240 >> minimums
print min_44080_82040 >> minimums
print min_44080_84840 >> minimums
print min_44080_87640 >> minimums
print min_44460_40040 >> minimums
print min_44460_42840 >> minimums
print min_44460_45640 >> minimums
print min_44460_48440 >> minimums
print min_44460_51240 >> minimums
print min_44460_54040 >> minimums
print min_44460_56840 >> minimums
print min_44460_59640 >> minimums
print min_44460_62440 >> minimums
print min_44460_65240 >> minimums
print min_44460_68040 >> minimums
print min_44460_70840 >> minimums
print min_44460_73640 >> minimums
print min_44460_76440 >> minimums
print min_44460_79240 >> minimums
print min_44460_82040 >> minimums
print min_44460_84840 >> minimums
print min_44460_87640 >> minimums
print min_44840_40040 >> minimums
print min_44840_42840 >> minimums
print min_44840_45640 >> minimums
print min_44840_48440 >> minimums
print min_44840_51240 >> minimums
print min_44840_54040 >> minimums
print min_44840_56840 >> minimums
print min_44840_59640 >> minimums
print min_44840_62440 >> minimums
print min_44840_65240 >> minimums
print min_44840_68040 >> minimums
print min_44840_70840 >> minimums
print min_44840_73640 >> minimums
print min_44840_76440 >> minimums
print min_44840_79240 >> minimums
print min_44840_82040 >> minimums
print min_44840_84840 >> minimums
print min_44840_87640 >> minimums
print min_45220_40040 >> minimums
print min_45220_42840 >> minimums
print min_45220_45640 >> minimums
print min_45220_48440 >> minimums
print min_45220_51240 >> minimums
print min_45220_54040 >> minimums
print min_45220_56840 >> minimums
print min_45220_59640 >> minimums
print min_45220_62440 >> minimums
print min_45220_65240 >> minimums
print min_45220_68040 >> minimums
print min_45220_70840 >> minimums
print min_45220_73640 >> minimums
print min_45220_76440 >> minimums
print min_45220_79240 >> minimums
print min_45220_82040 >> minimums
print min_45220_84840 >> minimums
print min_45220_87640 >> minimums
print min_45600_40040 >> minimums
print min_45600_42840 >> minimums
print min_45600_45640 >> minimums
print min_45600_48440 >> minimums
print min_45600_51240 >> minimums
print min_45600_54040 >> minimums
print min_45600_56840 >> minimums
print min_45600_59640 >> minimums
print min_45600_62440 >> minimums
print min_45600_65240 >> minimums
print min_45600_68040 >> minimums
print min_45600_70840 >> minimums
print min_45600_73640 >> minimums
print min_45600_76440 >> minimums
print min_45600_79240 >> minimums
print min_45600_82040 >> minimums
print min_45600_84840 >> minimums
print min_45600_87640 >> minimums
print min_46360_40040 >> minimums
print min_46360_42840 >> minimums
print min_46360_45640 >> minimums
print min_46360_48440 >> minimums
print min_46360_51240 >> minimums
print min_46360_54040 >> minimums
print min_46360_56840 >> minimums
print min_46360_59640 >> minimums
print min_46360_62440 >> minimums
print min_46360_65240 >> minimums
print min_46360_68040 >> minimums
print min_46360_70840 >> minimums
print min_46360_73640 >> minimums
print min_46360_76440 >> minimums
print min_46360_79240 >> minimums
print min_46360_82040 >> minimums
print min_46360_84840 >> minimums
print min_46360_87640 >> minimums
print min_46740_40040 >> minimums
print min_46740_42840 >> minimums
print min_46740_45640 >> minimums
print min_46740_48440 >> minimums
print min_46740_51240 >> minimums
print min_46740_54040 >> minimums
print min_46740_56840 >> minimums
print min_46740_59640 >> minimums
print min_46740_62440 >> minimums
print min_46740_65240 >> minimums
print min_46740_68040 >> minimums
print min_46740_70840 >> minimums
print min_46740_73640 >> minimums
print min_46740_76440 >> minimums
print min_46740_79240 >> minimums
print min_46740_82040 >> minimums
print min_46740_84840 >> minimums
print min_46740_87640 >> minimums
print min_47120_40040 >> minimums
print min_47120_42840 >> minimums
print min_47120_45640 >> minimums
print min_47120_48440 >> minimums
print min_47120_51240 >> minimums
print min_47120_54040 >> minimums
print min_47120_56840 >> minimums
print min_47120_59640 >> minimums
print min_47120_62440 >> minimums
print min_47120_65240 >> minimums
print min_47120_68040 >> minimums
print min_47120_70840 >> minimums
print min_47120_73640 >> minimums
print min_47120_76440 >> minimums
print min_47120_79240 >> minimums
print min_47120_82040 >> minimums
print min_47120_84840 >> minimums
print min_47120_87640 >> minimums
print min_47500_40040 >> minimums
print min_47500_42840 >> minimums
print min_47500_45640 >> minimums
print min_47500_48440 >> minimums
print min_47500_51240 >> minimums
print min_47500_54040 >> minimums
print min_47500_56840 >> minimums
print min_47500_59640 >> minimums
print min_47500_62440 >> minimums
print min_47500_65240 >> minimums
print min_47500_68040 >> minimums
print min_47500_70840 >> minimums
print min_47500_73640 >> minimums
print min_47500_76440 >> minimums
print min_47500_79240 >> minimums
print min_47500_82040 >> minimums
print min_47500_84840 >> minimums
print min_47500_87640 >> minimums
print min_47880_40040 >> minimums
print min_47880_42840 >> minimums
print min_47880_45640 >> minimums
print min_47880_48440 >> minimums
print min_47880_51240 >> minimums
print min_47880_54040 >> minimums
print min_47880_56840 >> minimums
print min_47880_59640 >> minimums
print min_47880_62440 >> minimums
print min_47880_65240 >> minimums
print min_47880_68040 >> minimums
print min_47880_70840 >> minimums
print min_47880_73640 >> minimums
print min_47880_76440 >> minimums
print min_47880_79240 >> minimums
print min_47880_82040 >> minimums
print min_47880_84840 >> minimums
print min_47880_87640 >> minimums
print min_48260_40040 >> minimums
print min_48260_42840 >> minimums
print min_48260_45640 >> minimums
print min_48260_48440 >> minimums
print min_48260_51240 >> minimums
print min_48260_54040 >> minimums
print min_48260_56840 >> minimums
print min_48260_59640 >> minimums
print min_48260_62440 >> minimums
print min_48260_65240 >> minimums
print min_48260_68040 >> minimums
print min_48260_70840 >> minimums
print min_48260_73640 >> minimums
print min_48260_76440 >> minimums
print min_48260_79240 >> minimums
print min_48260_82040 >> minimums
print min_48260_84840 >> minimums
print min_48260_87640 >> minimums
print min_48640_40040 >> minimums
print min_48640_42840 >> minimums
print min_48640_45640 >> minimums
print min_48640_48440 >> minimums
print min_48640_51240 >> minimums
print min_48640_54040 >> minimums
print min_48640_56840 >> minimums
print min_48640_59640 >> minimums
print min_48640_62440 >> minimums
print min_48640_65240 >> minimums
print min_48640_68040 >> minimums
print min_48640_70840 >> minimums
print min_48640_73640 >> minimums
print min_48640_76440 >> minimums
print min_48640_79240 >> minimums
print min_48640_82040 >> minimums
print min_48640_84840 >> minimums
print min_48640_87640 >> minimums
print min_49020_40040 >> minimums
print min_49020_42840 >> minimums
print min_49020_45640 >> minimums
print min_49020_48440 >> minimums
print min_49020_51240 >> minimums
print min_49020_54040 >> minimums
print min_49020_56840 >> minimums
print min_49020_59640 >> minimums
print min_49020_62440 >> minimums
print min_49020_65240 >> minimums
print min_49020_68040 >> minimums
print min_49020_70840 >> minimums
print min_49020_73640 >> minimums
print min_49020_76440 >> minimums
print min_49020_79240 >> minimums
print min_49020_82040 >> minimums
print min_49020_84840 >> minimums
print min_49020_87640 >> minimums
print min_49400_40040 >> minimums
print min_49400_42840 >> minimums
print min_49400_45640 >> minimums
print min_49400_48440 >> minimums
print min_49400_51240 >> minimums
print min_49400_54040 >> minimums
print min_49400_56840 >> minimums
print min_49400_59640 >> minimums
print min_49400_62440 >> minimums
print min_49400_65240 >> minimums
print min_49400_68040 >> minimums
print min_49400_70840 >> minimums
print min_49400_73640 >> minimums
print min_49400_76440 >> minimums
print min_49400_79240 >> minimums
print min_49400_82040 >> minimums
print min_49400_84840 >> minimums
print min_49400_87640 >> minimums
print min_49780_40040 >> minimums
print min_49780_42840 >> minimums
print min_49780_45640 >> minimums
print min_49780_48440 >> minimums
print min_49780_51240 >> minimums
print min_49780_54040 >> minimums
print min_49780_56840 >> minimums
print min_49780_59640 >> minimums
print min_49780_62440 >> minimums
print min_49780_65240 >> minimums
print min_49780_68040 >> minimums
print min_49780_70840 >> minimums
print min_49780_73640 >> minimums
print min_49780_76440 >> minimums
print min_49780_79240 >> minimums
print min_49780_82040 >> minimums
print min_49780_84840 >> minimums
print min_49780_87640 >> minimums
print min_50160_40040 >> minimums
print min_50160_42840 >> minimums
print min_50160_45640 >> minimums
print min_50160_48440 >> minimums
print min_50160_51240 >> minimums
print min_50160_54040 >> minimums
print min_50160_56840 >> minimums
print min_50160_59640 >> minimums
print min_50160_62440 >> minimums
print min_50160_65240 >> minimums
print min_50160_68040 >> minimums
print min_50160_70840 >> minimums
print min_50160_73640 >> minimums
print min_50160_76440 >> minimums
print min_50160_79240 >> minimums
print min_50160_82040 >> minimums
print min_50160_84840 >> minimums
print min_50160_87640 >> minimums
print min_50540_40040 >> minimums
print min_50540_42840 >> minimums
print min_50540_45640 >> minimums
print min_50540_48440 >> minimums
print min_50540_51240 >> minimums
print min_50540_54040 >> minimums
print min_50540_56840 >> minimums
print min_50540_59640 >> minimums
print min_50540_62440 >> minimums
print min_50540_65240 >> minimums
print min_50540_68040 >> minimums
print min_50540_70840 >> minimums
print min_50540_73640 >> minimums
print min_50540_76440 >> minimums
print min_50540_79240 >> minimums
print min_50540_82040 >> minimums
print min_50540_84840 >> minimums
print min_50540_87640 >> minimums
print min_50920_40040 >> minimums
print min_50920_42840 >> minimums
print min_50920_45640 >> minimums
print min_50920_48440 >> minimums
print min_50920_51240 >> minimums
print min_50920_54040 >> minimums
print min_50920_56840 >> minimums
print min_50920_59640 >> minimums
print min_50920_62440 >> minimums
print min_50920_65240 >> minimums
print min_50920_68040 >> minimums
print min_50920_70840 >> minimums
print min_50920_73640 >> minimums
print min_50920_76440 >> minimums
print min_50920_79240 >> minimums
print min_50920_82040 >> minimums
print min_50920_84840 >> minimums
print min_50920_87640 >> minimums
print min_51300_40040 >> minimums
print min_51300_42840 >> minimums
print min_51300_45640 >> minimums
print min_51300_48440 >> minimums
print min_51300_51240 >> minimums
print min_51300_54040 >> minimums
print min_51300_56840 >> minimums
print min_51300_59640 >> minimums
print min_51300_62440 >> minimums
print min_51300_65240 >> minimums
print min_51300_68040 >> minimums
print min_51300_70840 >> minimums
print min_51300_73640 >> minimums
print min_51300_76440 >> minimums
print min_51300_79240 >> minimums
print min_51300_82040 >> minimums
print min_51300_84840 >> minimums
print min_51300_87640 >> minimums
print min_51680_40040 >> minimums
print min_51680_42840 >> minimums
print min_51680_45640 >> minimums
print min_51680_48440 >> minimums
print min_51680_51240 >> minimums
print min_51680_54040 >> minimums
print min_51680_56840 >> minimums
print min_51680_59640 >> minimums
print min_51680_62440 >> minimums
print min_51680_65240 >> minimums
print min_51680_68040 >> minimums
print min_51680_70840 >> minimums
print min_51680_73640 >> minimums
print min_51680_76440 >> minimums
print min_51680_79240 >> minimums
print min_51680_82040 >> minimums
print min_51680_84840 >> minimums
print min_51680_87640 >> minimums
print min_52060_40040 >> minimums
print min_52060_42840 >> minimums
print min_52060_45640 >> minimums
print min_52060_48440 >> minimums
print min_52060_51240 >> minimums
print min_52060_54040 >> minimums
print min_52060_56840 >> minimums
print min_52060_59640 >> minimums
print min_52060_62440 >> minimums
print min_52060_65240 >> minimums
print min_52060_68040 >> minimums
print min_52060_70840 >> minimums
print min_52060_73640 >> minimums
print min_52060_76440 >> minimums
print min_52060_79240 >> minimums
print min_52060_82040 >> minimums
print min_52060_84840 >> minimums
print min_52060_87640 >> minimums
print min_52440_40040 >> minimums
print min_52440_42840 >> minimums
print min_52440_45640 >> minimums
print min_52440_48440 >> minimums
print min_52440_51240 >> minimums
print min_52440_54040 >> minimums
print min_52440_56840 >> minimums
print min_52440_59640 >> minimums
print min_52440_62440 >> minimums
print min_52440_65240 >> minimums
print min_52440_68040 >> minimums
print min_52440_70840 >> minimums
print min_52440_73640 >> minimums
print min_52440_76440 >> minimums
print min_52440_79240 >> minimums
print min_52440_82040 >> minimums
print min_52440_84840 >> minimums
print min_52440_87640 >> minimums
print min_52820_40040 >> minimums
print min_52820_42840 >> minimums
print min_52820_45640 >> minimums
print min_52820_48440 >> minimums
print min_52820_51240 >> minimums
print min_52820_54040 >> minimums
print min_52820_56840 >> minimums
print min_52820_59640 >> minimums
print min_52820_62440 >> minimums
print min_52820_65240 >> minimums
print min_52820_68040 >> minimums
print min_52820_70840 >> minimums
print min_52820_73640 >> minimums
print min_52820_76440 >> minimums
print min_52820_79240 >> minimums
print min_52820_82040 >> minimums
print min_52820_84840 >> minimums
print min_52820_87640 >> minimums
print min_53200_40040 >> minimums
print min_53200_42840 >> minimums
print min_53200_45640 >> minimums
print min_53200_48440 >> minimums
print min_53200_51240 >> minimums
print min_53200_54040 >> minimums
print min_53200_56840 >> minimums
print min_53200_59640 >> minimums
print min_53200_62440 >> minimums
print min_53200_65240 >> minimums
print min_53200_68040 >> minimums
print min_53200_70840 >> minimums
print min_53200_73640 >> minimums
print min_53200_76440 >> minimums
print min_53200_79240 >> minimums
print min_53200_82040 >> minimums
print min_53200_84840 >> minimums
print min_53200_87640 >> minimums
print min_53580_40040 >> minimums
print min_53580_42840 >> minimums
print min_53580_45640 >> minimums
print min_53580_48440 >> minimums
print min_53580_51240 >> minimums
print min_53580_54040 >> minimums
print min_53580_56840 >> minimums
print min_53580_59640 >> minimums
print min_53580_62440 >> minimums
print min_53580_65240 >> minimums
print min_53580_68040 >> minimums
print min_53580_70840 >> minimums
print min_53580_73640 >> minimums
print min_53580_76440 >> minimums
print min_53580_79240 >> minimums
print min_53580_82040 >> minimums
print min_53580_84840 >> minimums
print min_53580_87640 >> minimums
print min_53960_40040 >> minimums
print min_53960_42840 >> minimums
print min_53960_45640 >> minimums
print min_53960_48440 >> minimums
print min_53960_51240 >> minimums
print min_53960_54040 >> minimums
print min_53960_56840 >> minimums
print min_53960_59640 >> minimums
print min_53960_62440 >> minimums
print min_53960_65240 >> minimums
print min_53960_68040 >> minimums
print min_53960_70840 >> minimums
print min_53960_73640 >> minimums
print min_53960_76440 >> minimums
print min_53960_79240 >> minimums
print min_53960_82040 >> minimums
print min_53960_84840 >> minimums
print min_53960_87640 >> minimums
print min_54340_40040 >> minimums
print min_54340_42840 >> minimums
print min_54340_45640 >> minimums
print min_54340_48440 >> minimums
print min_54340_51240 >> minimums
print min_54340_54040 >> minimums
print min_54340_56840 >> minimums
print min_54340_59640 >> minimums
print min_54340_62440 >> minimums
print min_54340_65240 >> minimums
print min_54340_68040 >> minimums
print min_54340_70840 >> minimums
print min_54340_73640 >> minimums
print min_54340_76440 >> minimums
print min_54340_79240 >> minimums
print min_54340_82040 >> minimums
print min_54340_84840 >> minimums
print min_54340_87640 >> minimums
print min_54720_40040 >> minimums
print min_54720_42840 >> minimums
print min_54720_45640 >> minimums
print min_54720_48440 >> minimums
print min_54720_51240 >> minimums
print min_54720_54040 >> minimums
print min_54720_56840 >> minimums
print min_54720_59640 >> minimums
print min_54720_62440 >> minimums
print min_54720_65240 >> minimums
print min_54720_68040 >> minimums
print min_54720_70840 >> minimums
print min_54720_73640 >> minimums
print min_54720_76440 >> minimums
print min_54720_79240 >> minimums
print min_54720_82040 >> minimums
print min_54720_84840 >> minimums
print min_54720_87640 >> minimums
print min_55100_40040 >> minimums
print min_55100_42840 >> minimums
print min_55100_45640 >> minimums
print min_55100_48440 >> minimums
print min_55100_51240 >> minimums
print min_55100_54040 >> minimums
print min_55100_56840 >> minimums
print min_55100_59640 >> minimums
print min_55100_62440 >> minimums
print min_55100_65240 >> minimums
print min_55100_68040 >> minimums
print min_55100_70840 >> minimums
print min_55100_73640 >> minimums
print min_55100_76440 >> minimums
print min_55100_79240 >> minimums
print min_55100_82040 >> minimums
print min_55100_84840 >> minimums
print min_55100_87640 >> minimums
print min_55480_40040 >> minimums
print min_55480_42840 >> minimums
print min_55480_45640 >> minimums
print min_55480_48440 >> minimums
print min_55480_51240 >> minimums
print min_55480_54040 >> minimums
print min_55480_56840 >> minimums
print min_55480_59640 >> minimums
print min_55480_62440 >> minimums
print min_55480_65240 >> minimums
print min_55480_68040 >> minimums
print min_55480_70840 >> minimums
print min_55480_73640 >> minimums
print min_55480_76440 >> minimums
print min_55480_79240 >> minimums
print min_55480_82040 >> minimums
print min_55480_84840 >> minimums
print min_55480_87640 >> minimums
print min_55860_40040 >> minimums
print min_55860_42840 >> minimums
print min_55860_45640 >> minimums
print min_55860_48440 >> minimums
print min_55860_51240 >> minimums
print min_55860_54040 >> minimums
print min_55860_56840 >> minimums
print min_55860_59640 >> minimums
print min_55860_62440 >> minimums
print min_55860_65240 >> minimums
print min_55860_68040 >> minimums
print min_55860_70840 >> minimums
print min_55860_73640 >> minimums
print min_55860_76440 >> minimums
print min_55860_79240 >> minimums
print min_55860_82040 >> minimums
print min_55860_84840 >> minimums
print min_55860_87640 >> minimums
print min_56240_40040 >> minimums
print min_56240_42840 >> minimums
print min_56240_45640 >> minimums
print min_56240_48440 >> minimums
print min_56240_51240 >> minimums
print min_56240_54040 >> minimums
print min_56240_56840 >> minimums
print min_56240_59640 >> minimums
print min_56240_62440 >> minimums
print min_56240_65240 >> minimums
print min_56240_68040 >> minimums
print min_56240_70840 >> minimums
print min_56240_73640 >> minimums
print min_56240_76440 >> minimums
print min_56240_79240 >> minimums
print min_56240_82040 >> minimums
print min_56240_84840 >> minimums
print min_56240_87640 >> minimums
print min_56620_40040 >> minimums
print min_56620_42840 >> minimums
print min_56620_45640 >> minimums
print min_56620_48440 >> minimums
print min_56620_51240 >> minimums
print min_56620_54040 >> minimums
print min_56620_56840 >> minimums
print min_56620_59640 >> minimums
print min_56620_62440 >> minimums
print min_56620_65240 >> minimums
print min_56620_68040 >> minimums
print min_56620_70840 >> minimums
print min_56620_73640 >> minimums
print min_56620_76440 >> minimums
print min_56620_79240 >> minimums
print min_56620_82040 >> minimums
print min_56620_84840 >> minimums
print min_56620_87640 >> minimums
print min_57000_40040 >> minimums
print min_57000_42840 >> minimums
print min_57000_45640 >> minimums
print min_57000_48440 >> minimums
print min_57000_51240 >> minimums
print min_57000_54040 >> minimums
print min_57000_56840 >> minimums
print min_57000_59640 >> minimums
print min_57000_62440 >> minimums
print min_57000_65240 >> minimums
print min_57000_68040 >> minimums
print min_57000_70840 >> minimums
print min_57000_73640 >> minimums
print min_57000_76440 >> minimums
print min_57000_79240 >> minimums
print min_57000_82040 >> minimums
print min_57000_84840 >> minimums
print min_57000_87640 >> minimums
print min_57380_40040 >> minimums
print min_57380_42840 >> minimums
print min_57380_45640 >> minimums
print min_57380_48440 >> minimums
print min_57380_51240 >> minimums
print min_57380_54040 >> minimums
print min_57380_56840 >> minimums
print min_57380_59640 >> minimums
print min_57380_62440 >> minimums
print min_57380_65240 >> minimums
print min_57380_68040 >> minimums
print min_57380_70840 >> minimums
print min_57380_73640 >> minimums
print min_57380_76440 >> minimums
print min_57380_79240 >> minimums
print min_57380_82040 >> minimums
print min_57380_84840 >> minimums
print min_57380_87640 >> minimums
print min_57760_40040 >> minimums
print min_57760_42840 >> minimums
print min_57760_45640 >> minimums
print min_57760_48440 >> minimums
print min_57760_51240 >> minimums
print min_57760_54040 >> minimums
print min_57760_56840 >> minimums
print min_57760_59640 >> minimums
print min_57760_62440 >> minimums
print min_57760_65240 >> minimums
print min_57760_68040 >> minimums
print min_57760_70840 >> minimums
print min_57760_73640 >> minimums
print min_57760_76440 >> minimums
print min_57760_79240 >> minimums
print min_57760_82040 >> minimums
print min_57760_84840 >> minimums
print min_57760_87640 >> minimums
print min_58140_40040 >> minimums
print min_58140_42840 >> minimums
print min_58140_45640 >> minimums
print min_58140_48440 >> minimums
print min_58140_51240 >> minimums
print min_58140_54040 >> minimums
print min_58140_56840 >> minimums
print min_58140_59640 >> minimums
print min_58140_62440 >> minimums
print min_58140_65240 >> minimums
print min_58140_68040 >> minimums
print min_58140_70840 >> minimums
print min_58140_73640 >> minimums
print min_58140_76440 >> minimums
print min_58140_79240 >> minimums
print min_58140_82040 >> minimums
print min_58140_84840 >> minimums
print min_58140_87640 >> minimums
print min_58520_40040 >> minimums
print min_58520_42840 >> minimums
print min_58520_45640 >> minimums
print min_58520_48440 >> minimums
print min_58520_51240 >> minimums
print min_58520_54040 >> minimums
print min_58520_56840 >> minimums
print min_58520_59640 >> minimums
print min_58520_62440 >> minimums
print min_58520_65240 >> minimums
print min_58520_68040 >> minimums
print min_58520_70840 >> minimums
print min_58520_73640 >> minimums
print min_58520_76440 >> minimums
print min_58520_79240 >> minimums
print min_58520_82040 >> minimums
print min_58520_84840 >> minimums
print min_58520_87640 >> minimums
print min_58900_40040 >> minimums
print min_58900_42840 >> minimums
print min_58900_45640 >> minimums
print min_58900_48440 >> minimums
print min_58900_51240 >> minimums
print min_58900_54040 >> minimums
print min_58900_56840 >> minimums
print min_58900_59640 >> minimums
print min_58900_62440 >> minimums
print min_58900_65240 >> minimums
print min_58900_68040 >> minimums
print min_58900_70840 >> minimums
print min_58900_73640 >> minimums
print min_58900_76440 >> minimums
print min_58900_79240 >> minimums
print min_58900_82040 >> minimums
print min_58900_84840 >> minimums
print min_58900_87640 >> minimums
print min_59280_40040 >> minimums
print min_59280_42840 >> minimums
print min_59280_45640 >> minimums
print min_59280_48440 >> minimums
print min_59280_51240 >> minimums
print min_59280_54040 >> minimums
print min_59280_56840 >> minimums
print min_59280_59640 >> minimums
print min_59280_62440 >> minimums
print min_59280_65240 >> minimums
print min_59280_68040 >> minimums
print min_59280_70840 >> minimums
print min_59280_73640 >> minimums
print min_59280_76440 >> minimums
print min_59280_79240 >> minimums
print min_59280_82040 >> minimums
print min_59280_84840 >> minimums
print min_59280_87640 >> minimums
print min_59660_40040 >> minimums
print min_59660_42840 >> minimums
print min_59660_45640 >> minimums
print min_59660_48440 >> minimums
print min_59660_51240 >> minimums
print min_59660_54040 >> minimums
print min_59660_56840 >> minimums
print min_59660_59640 >> minimums
print min_59660_62440 >> minimums
print min_59660_65240 >> minimums
print min_59660_68040 >> minimums
print min_59660_70840 >> minimums
print min_59660_73640 >> minimums
print min_59660_76440 >> minimums
print min_59660_79240 >> minimums
print min_59660_82040 >> minimums
print min_59660_84840 >> minimums
print min_59660_87640 >> minimums
print min_60040_40040 >> minimums
print min_60040_42840 >> minimums
print min_60040_45640 >> minimums
print min_60040_48440 >> minimums
print min_60040_51240 >> minimums
print min_60040_54040 >> minimums
print min_60040_56840 >> minimums
print min_60040_59640 >> minimums
print min_60040_62440 >> minimums
print min_60040_65240 >> minimums
print min_60040_68040 >> minimums
print min_60040_70840 >> minimums
print min_60040_73640 >> minimums
print min_60040_76440 >> minimums
print min_60040_79240 >> minimums
print min_60040_82040 >> minimums
print min_60040_84840 >> minimums
print min_60040_87640 >> minimums
print min_60420_40040 >> minimums
print min_60420_42840 >> minimums
print min_60420_45640 >> minimums
print min_60420_48440 >> minimums
print min_60420_51240 >> minimums
print min_60420_54040 >> minimums
print min_60420_56840 >> minimums
print min_60420_59640 >> minimums
print min_60420_62440 >> minimums
print min_60420_65240 >> minimums
print min_60420_68040 >> minimums
print min_60420_70840 >> minimums
print min_60420_73640 >> minimums
print min_60420_76440 >> minimums
print min_60420_79240 >> minimums
print min_60420_82040 >> minimums
print min_60420_84840 >> minimums
print min_60420_87640 >> minimums
print min_60800_40040 >> minimums
print min_60800_42840 >> minimums
print min_60800_45640 >> minimums
print min_60800_48440 >> minimums
print min_60800_51240 >> minimums
print min_60800_54040 >> minimums
print min_60800_56840 >> minimums
print min_60800_59640 >> minimums
print min_60800_62440 >> minimums
print min_60800_65240 >> minimums
print min_60800_68040 >> minimums
print min_60800_70840 >> minimums
print min_60800_73640 >> minimums
print min_60800_76440 >> minimums
print min_60800_79240 >> minimums
print min_60800_82040 >> minimums
print min_60800_84840 >> minimums
print min_60800_87640 >> minimums
print min_61180_40040 >> minimums
print min_61180_42840 >> minimums
print min_61180_45640 >> minimums
print min_61180_48440 >> minimums
print min_61180_51240 >> minimums
print min_61180_54040 >> minimums
print min_61180_56840 >> minimums
print min_61180_59640 >> minimums
print min_61180_62440 >> minimums
print min_61180_65240 >> minimums
print min_61180_68040 >> minimums
print min_61180_70840 >> minimums
print min_61180_73640 >> minimums
print min_61180_76440 >> minimums
print min_61180_79240 >> minimums
print min_61180_82040 >> minimums
print min_61180_84840 >> minimums
print min_61180_87640 >> minimums
print min_61560_40040 >> minimums
print min_61560_42840 >> minimums
print min_61560_45640 >> minimums
print min_61560_48440 >> minimums
print min_61560_51240 >> minimums
print min_61560_54040 >> minimums
print min_61560_56840 >> minimums
print min_61560_59640 >> minimums
print min_61560_62440 >> minimums
print min_61560_65240 >> minimums
print min_61560_68040 >> minimums
print min_61560_70840 >> minimums
print min_61560_73640 >> minimums
print min_61560_76440 >> minimums
print min_61560_79240 >> minimums
print min_61560_82040 >> minimums
print min_61560_84840 >> minimums
print min_61560_87640 >> minimums
print min_61940_40040 >> minimums
print min_61940_42840 >> minimums
print min_61940_45640 >> minimums
print min_61940_48440 >> minimums
print min_61940_51240 >> minimums
print min_61940_54040 >> minimums
print min_61940_56840 >> minimums
print min_61940_59640 >> minimums
print min_61940_62440 >> minimums
print min_61940_65240 >> minimums
print min_61940_68040 >> minimums
print min_61940_70840 >> minimums
print min_61940_73640 >> minimums
print min_61940_76440 >> minimums
print min_61940_79240 >> minimums
print min_61940_82040 >> minimums
print min_61940_84840 >> minimums
print min_61940_87640 >> minimums
print min_62320_40040 >> minimums
print min_62320_42840 >> minimums
print min_62320_45640 >> minimums
print min_62320_48440 >> minimums
print min_62320_51240 >> minimums
print min_62320_54040 >> minimums
print min_62320_56840 >> minimums
print min_62320_59640 >> minimums
print min_62320_62440 >> minimums
print min_62320_65240 >> minimums
print min_62320_68040 >> minimums
print min_62320_70840 >> minimums
print min_62320_73640 >> minimums
print min_62320_76440 >> minimums
print min_62320_79240 >> minimums
print min_62320_82040 >> minimums
print min_62320_84840 >> minimums
print min_62320_87640 >> minimums
print min_63080_40040 >> minimums
print min_63080_42840 >> minimums
print min_63080_45640 >> minimums
print min_63080_48440 >> minimums
print min_63080_51240 >> minimums
print min_63080_54040 >> minimums
print min_63080_56840 >> minimums
print min_63080_59640 >> minimums
print min_63080_62440 >> minimums
print min_63080_65240 >> minimums
print min_63080_68040 >> minimums
print min_63080_70840 >> minimums
print min_63080_73640 >> minimums
print min_63080_76440 >> minimums
print min_63080_79240 >> minimums
print min_63080_82040 >> minimums
print min_63080_84840 >> minimums
print min_63080_87640 >> minimums
print min_63460_40040 >> minimums
print min_63460_42840 >> minimums
print min_63460_45640 >> minimums
print min_63460_48440 >> minimums
print min_63460_51240 >> minimums
print min_63460_54040 >> minimums
print min_63460_56840 >> minimums
print min_63460_59640 >> minimums
print min_63460_62440 >> minimums
print min_63460_65240 >> minimums
print min_63460_68040 >> minimums
print min_63460_70840 >> minimums
print min_63460_73640 >> minimums
print min_63460_76440 >> minimums
print min_63460_79240 >> minimums
print min_63460_82040 >> minimums
print min_63460_84840 >> minimums
print min_63460_87640 >> minimums
print min_63840_40040 >> minimums
print min_63840_42840 >> minimums
print min_63840_45640 >> minimums
print min_63840_48440 >> minimums
print min_63840_51240 >> minimums
print min_63840_54040 >> minimums
print min_63840_56840 >> minimums
print min_63840_59640 >> minimums
print min_63840_62440 >> minimums
print min_63840_65240 >> minimums
print min_63840_68040 >> minimums
print min_63840_70840 >> minimums
print min_63840_73640 >> minimums
print min_63840_76440 >> minimums
print min_63840_79240 >> minimums
print min_63840_82040 >> minimums
print min_63840_84840 >> minimums
print min_63840_87640 >> minimums
print min_64220_40040 >> minimums
print min_64220_42840 >> minimums
print min_64220_45640 >> minimums
print min_64220_48440 >> minimums
print min_64220_51240 >> minimums
print min_64220_54040 >> minimums
print min_64220_56840 >> minimums
print min_64220_59640 >> minimums
print min_64220_62440 >> minimums
print min_64220_65240 >> minimums
print min_64220_68040 >> minimums
print min_64220_70840 >> minimums
print min_64220_73640 >> minimums
print min_64220_76440 >> minimums
print min_64220_79240 >> minimums
print min_64220_82040 >> minimums
print min_64220_84840 >> minimums
print min_64220_87640 >> minimums
print min_64600_40040 >> minimums
print min_64600_42840 >> minimums
print min_64600_45640 >> minimums
print min_64600_48440 >> minimums
print min_64600_51240 >> minimums
print min_64600_54040 >> minimums
print min_64600_56840 >> minimums
print min_64600_59640 >> minimums
print min_64600_62440 >> minimums
print min_64600_65240 >> minimums
print min_64600_68040 >> minimums
print min_64600_70840 >> minimums
print min_64600_73640 >> minimums
print min_64600_76440 >> minimums
print min_64600_79240 >> minimums
print min_64600_82040 >> minimums
print min_64600_84840 >> minimums
print min_64600_87640 >> minimums
print min_64980_40040 >> minimums
print min_64980_42840 >> minimums
print min_64980_45640 >> minimums
print min_64980_48440 >> minimums
print min_64980_51240 >> minimums
print min_64980_54040 >> minimums
print min_64980_56840 >> minimums
print min_64980_59640 >> minimums
print min_64980_62440 >> minimums
print min_64980_65240 >> minimums
print min_64980_68040 >> minimums
print min_64980_70840 >> minimums
print min_64980_73640 >> minimums
print min_64980_76440 >> minimums
print min_64980_79240 >> minimums
print min_64980_82040 >> minimums
print min_64980_84840 >> minimums
print min_64980_87640 >> minimums
print min_65360_40040 >> minimums
print min_65360_42840 >> minimums
print min_65360_45640 >> minimums
print min_65360_48440 >> minimums
print min_65360_51240 >> minimums
print min_65360_54040 >> minimums
print min_65360_56840 >> minimums
print min_65360_59640 >> minimums
print min_65360_62440 >> minimums
print min_65360_65240 >> minimums
print min_65360_68040 >> minimums
print min_65360_70840 >> minimums
print min_65360_73640 >> minimums
print min_65360_76440 >> minimums
print min_65360_79240 >> minimums
print min_65360_82040 >> minimums
print min_65360_84840 >> minimums
print min_65360_87640 >> minimums
print min_65740_40040 >> minimums
print min_65740_42840 >> minimums
print min_65740_45640 >> minimums
print min_65740_48440 >> minimums
print min_65740_51240 >> minimums
print min_65740_54040 >> minimums
print min_65740_56840 >> minimums
print min_65740_59640 >> minimums
print min_65740_62440 >> minimums
print min_65740_65240 >> minimums
print min_65740_68040 >> minimums
print min_65740_70840 >> minimums
print min_65740_73640 >> minimums
print min_65740_76440 >> minimums
print min_65740_79240 >> minimums
print min_65740_82040 >> minimums
print min_65740_84840 >> minimums
print min_65740_87640 >> minimums
print min_66120_40040 >> minimums
print min_66120_42840 >> minimums
print min_66120_45640 >> minimums
print min_66120_48440 >> minimums
print min_66120_51240 >> minimums
print min_66120_54040 >> minimums
print min_66120_56840 >> minimums
print min_66120_59640 >> minimums
print min_66120_62440 >> minimums
print min_66120_65240 >> minimums
print min_66120_68040 >> minimums
print min_66120_70840 >> minimums
print min_66120_73640 >> minimums
print min_66120_76440 >> minimums
print min_66120_79240 >> minimums
print min_66120_82040 >> minimums
print min_66120_84840 >> minimums
print min_66120_87640 >> minimums
print min_66880_40040 >> minimums
print min_66880_42840 >> minimums
print min_66880_45640 >> minimums
print min_66880_48440 >> minimums
print min_66880_51240 >> minimums
print min_66880_54040 >> minimums
print min_66880_56840 >> minimums
print min_66880_59640 >> minimums
print min_66880_62440 >> minimums
print min_66880_65240 >> minimums
print min_66880_68040 >> minimums
print min_66880_70840 >> minimums
print min_66880_73640 >> minimums
print min_66880_76440 >> minimums
print min_66880_79240 >> minimums
print min_66880_82040 >> minimums
print min_66880_84840 >> minimums
print min_66880_87640 >> minimums
print min_67260_40040 >> minimums
print min_67260_42840 >> minimums
print min_67260_45640 >> minimums
print min_67260_48440 >> minimums
print min_67260_51240 >> minimums
print min_67260_54040 >> minimums
print min_67260_56840 >> minimums
print min_67260_59640 >> minimums
print min_67260_62440 >> minimums
print min_67260_65240 >> minimums
print min_67260_68040 >> minimums
print min_67260_70840 >> minimums
print min_67260_73640 >> minimums
print min_67260_76440 >> minimums
print min_67260_79240 >> minimums
print min_67260_82040 >> minimums
print min_67260_84840 >> minimums
print min_67260_87640 >> minimums
print min_68020_40040 >> minimums
print min_68020_42840 >> minimums
print min_68020_45640 >> minimums
print min_68020_48440 >> minimums
print min_68020_51240 >> minimums
print min_68020_54040 >> minimums
print min_68020_56840 >> minimums
print min_68020_59640 >> minimums
print min_68020_62440 >> minimums
print min_68020_65240 >> minimums
print min_68020_68040 >> minimums
print min_68020_70840 >> minimums
print min_68020_73640 >> minimums
print min_68020_76440 >> minimums
print min_68020_79240 >> minimums
print min_68020_82040 >> minimums
print min_68020_84840 >> minimums
print min_68020_87640 >> minimums
print min_68400_40040 >> minimums
print min_68400_42840 >> minimums
print min_68400_45640 >> minimums
print min_68400_48440 >> minimums
print min_68400_51240 >> minimums
print min_68400_54040 >> minimums
print min_68400_56840 >> minimums
print min_68400_59640 >> minimums
print min_68400_62440 >> minimums
print min_68400_65240 >> minimums
print min_68400_68040 >> minimums
print min_68400_70840 >> minimums
print min_68400_73640 >> minimums
print min_68400_76440 >> minimums
print min_68400_79240 >> minimums
print min_68400_82040 >> minimums
print min_68400_84840 >> minimums
print min_68400_87640 >> minimums
print min_68780_40040 >> minimums
print min_68780_42840 >> minimums
print min_68780_45640 >> minimums
print min_68780_48440 >> minimums
print min_68780_51240 >> minimums
print min_68780_54040 >> minimums
print min_68780_56840 >> minimums
print min_68780_59640 >> minimums
print min_68780_62440 >> minimums
print min_68780_65240 >> minimums
print min_68780_68040 >> minimums
print min_68780_70840 >> minimums
print min_68780_73640 >> minimums
print min_68780_76440 >> minimums
print min_68780_79240 >> minimums
print min_68780_82040 >> minimums
print min_68780_84840 >> minimums
print min_68780_87640 >> minimums
print min_69160_40040 >> minimums
print min_69160_42840 >> minimums
print min_69160_45640 >> minimums
print min_69160_48440 >> minimums
print min_69160_51240 >> minimums
print min_69160_54040 >> minimums
print min_69160_56840 >> minimums
print min_69160_59640 >> minimums
print min_69160_62440 >> minimums
print min_69160_65240 >> minimums
print min_69160_68040 >> minimums
print min_69160_70840 >> minimums
print min_69160_73640 >> minimums
print min_69160_76440 >> minimums
print min_69160_79240 >> minimums
print min_69160_82040 >> minimums
print min_69160_84840 >> minimums
print min_69160_87640 >> minimums
print min_69920_40040 >> minimums
print min_69920_42840 >> minimums
print min_69920_45640 >> minimums
print min_69920_48440 >> minimums
print min_69920_51240 >> minimums
print min_69920_54040 >> minimums
print min_69920_56840 >> minimums
print min_69920_59640 >> minimums
print min_69920_62440 >> minimums
print min_69920_65240 >> minimums
print min_69920_68040 >> minimums
print min_69920_70840 >> minimums
print min_69920_73640 >> minimums
print min_69920_76440 >> minimums
print min_69920_79240 >> minimums
print min_69920_82040 >> minimums
print min_69920_84840 >> minimums
print min_69920_87640 >> minimums
print min_70300_40040 >> minimums
print min_70300_42840 >> minimums
print min_70300_45640 >> minimums
print min_70300_48440 >> minimums
print min_70300_51240 >> minimums
print min_70300_54040 >> minimums
print min_70300_56840 >> minimums
print min_70300_59640 >> minimums
print min_70300_62440 >> minimums
print min_70300_65240 >> minimums
print min_70300_68040 >> minimums
print min_70300_70840 >> minimums
print min_70300_73640 >> minimums
print min_70300_76440 >> minimums
print min_70300_79240 >> minimums
print min_70300_82040 >> minimums
print min_70300_84840 >> minimums
print min_70300_87640 >> minimums
print min_71060_40040 >> minimums
print min_71060_42840 >> minimums
print min_71060_45640 >> minimums
print min_71060_48440 >> minimums
print min_71060_51240 >> minimums
print min_71060_54040 >> minimums
print min_71060_56840 >> minimums
print min_71060_59640 >> minimums
print min_71060_62440 >> minimums
print min_71060_65240 >> minimums
print min_71060_68040 >> minimums
print min_71060_70840 >> minimums
print min_71060_73640 >> minimums
print min_71060_76440 >> minimums
print min_71060_79240 >> minimums
print min_71060_82040 >> minimums
print min_71060_84840 >> minimums
print min_71060_87640 >> minimums
print min_71820_40040 >> minimums
print min_71820_42840 >> minimums
print min_71820_45640 >> minimums
print min_71820_48440 >> minimums
print min_71820_51240 >> minimums
print min_71820_54040 >> minimums
print min_71820_56840 >> minimums
print min_71820_59640 >> minimums
print min_71820_62440 >> minimums
print min_71820_65240 >> minimums
print min_71820_68040 >> minimums
print min_71820_70840 >> minimums
print min_71820_73640 >> minimums
print min_71820_76440 >> minimums
print min_71820_79240 >> minimums
print min_71820_82040 >> minimums
print min_71820_84840 >> minimums
print min_71820_87640 >> minimums
print min_72200_40040 >> minimums
print min_72200_42840 >> minimums
print min_72200_45640 >> minimums
print min_72200_48440 >> minimums
print min_72200_51240 >> minimums
print min_72200_54040 >> minimums
print min_72200_56840 >> minimums
print min_72200_59640 >> minimums
print min_72200_62440 >> minimums
print min_72200_65240 >> minimums
print min_72200_68040 >> minimums
print min_72200_70840 >> minimums
print min_72200_73640 >> minimums
print min_72200_76440 >> minimums
print min_72200_79240 >> minimums
print min_72200_82040 >> minimums
print min_72200_84840 >> minimums
print min_72200_87640 >> minimums
print min_72960_40040 >> minimums
print min_72960_42840 >> minimums
print min_72960_45640 >> minimums
print min_72960_48440 >> minimums
print min_72960_51240 >> minimums
print min_72960_54040 >> minimums
print min_72960_56840 >> minimums
print min_72960_59640 >> minimums
print min_72960_62440 >> minimums
print min_72960_65240 >> minimums
print min_72960_68040 >> minimums
print min_72960_70840 >> minimums
print min_72960_73640 >> minimums
print min_72960_76440 >> minimums
print min_72960_79240 >> minimums
print min_72960_82040 >> minimums
print min_72960_84840 >> minimums
print min_72960_87640 >> minimums
print min_73340_40040 >> minimums
print min_73340_42840 >> minimums
print min_73340_45640 >> minimums
print min_73340_48440 >> minimums
print min_73340_51240 >> minimums
print min_73340_54040 >> minimums
print min_73340_56840 >> minimums
print min_73340_59640 >> minimums
print min_73340_62440 >> minimums
print min_73340_65240 >> minimums
print min_73340_68040 >> minimums
print min_73340_70840 >> minimums
print min_73340_73640 >> minimums
print min_73340_76440 >> minimums
print min_73340_79240 >> minimums
print min_73340_82040 >> minimums
print min_73340_84840 >> minimums
print min_73340_87640 >> minimums
print min_73720_40040 >> minimums
print min_73720_42840 >> minimums
print min_73720_45640 >> minimums
print min_73720_48440 >> minimums
print min_73720_51240 >> minimums
print min_73720_54040 >> minimums
print min_73720_56840 >> minimums
print min_73720_59640 >> minimums
print min_73720_62440 >> minimums
print min_73720_65240 >> minimums
print min_73720_68040 >> minimums
print min_73720_70840 >> minimums
print min_73720_73640 >> minimums
print min_73720_76440 >> minimums
print min_73720_79240 >> minimums
print min_73720_82040 >> minimums
print min_73720_84840 >> minimums
print min_73720_87640 >> minimums
print min_74100_40040 >> minimums
print min_74100_42840 >> minimums
print min_74100_45640 >> minimums
print min_74100_48440 >> minimums
print min_74100_51240 >> minimums
print min_74100_54040 >> minimums
print min_74100_56840 >> minimums
print min_74100_59640 >> minimums
print min_74100_62440 >> minimums
print min_74100_65240 >> minimums
print min_74100_68040 >> minimums
print min_74100_70840 >> minimums
print min_74100_73640 >> minimums
print min_74100_76440 >> minimums
print min_74100_79240 >> minimums
print min_74100_82040 >> minimums
print min_74100_84840 >> minimums
print min_74100_87640 >> minimums
print min_74860_40040 >> minimums
print min_74860_42840 >> minimums
print min_74860_45640 >> minimums
print min_74860_48440 >> minimums
print min_74860_51240 >> minimums
print min_74860_54040 >> minimums
print min_74860_56840 >> minimums
print min_74860_59640 >> minimums
print min_74860_62440 >> minimums
print min_74860_65240 >> minimums
print min_74860_68040 >> minimums
print min_74860_70840 >> minimums
print min_74860_73640 >> minimums
print min_74860_76440 >> minimums
print min_74860_79240 >> minimums
print min_74860_82040 >> minimums
print min_74860_84840 >> minimums
print min_74860_87640 >> minimums
print min_75240_40040 >> minimums
print min_75240_42840 >> minimums
print min_75240_45640 >> minimums
print min_75240_48440 >> minimums
print min_75240_51240 >> minimums
print min_75240_54040 >> minimums
print min_75240_56840 >> minimums
print min_75240_59640 >> minimums
print min_75240_62440 >> minimums
print min_75240_65240 >> minimums
print min_75240_68040 >> minimums
print min_75240_70840 >> minimums
print min_75240_73640 >> minimums
print min_75240_76440 >> minimums
print min_75240_79240 >> minimums
print min_75240_82040 >> minimums
print min_75240_84840 >> minimums
print min_75240_87640 >> minimums
print min_76000_40040 >> minimums
print min_76000_42840 >> minimums
print min_76000_45640 >> minimums
print min_76000_48440 >> minimums
print min_76000_51240 >> minimums
print min_76000_54040 >> minimums
print min_76000_56840 >> minimums
print min_76000_59640 >> minimums
print min_76000_62440 >> minimums
print min_76000_65240 >> minimums
print min_76000_68040 >> minimums
print min_76000_70840 >> minimums
print min_76000_73640 >> minimums
print min_76000_76440 >> minimums
print min_76000_79240 >> minimums
print min_76000_82040 >> minimums
print min_76000_84840 >> minimums
print min_76000_87640 >> minimums
print min_76380_40040 >> minimums
print min_76380_42840 >> minimums
print min_76380_45640 >> minimums
print min_76380_48440 >> minimums
print min_76380_51240 >> minimums
print min_76380_54040 >> minimums
print min_76380_56840 >> minimums
print min_76380_59640 >> minimums
print min_76380_62440 >> minimums
print min_76380_65240 >> minimums
print min_76380_68040 >> minimums
print min_76380_70840 >> minimums
print min_76380_73640 >> minimums
print min_76380_76440 >> minimums
print min_76380_79240 >> minimums
print min_76380_82040 >> minimums
print min_76380_84840 >> minimums
print min_76380_87640 >> minimums
print min_76760_40040 >> minimums
print min_76760_42840 >> minimums
print min_76760_45640 >> minimums
print min_76760_48440 >> minimums
print min_76760_51240 >> minimums
print min_76760_54040 >> minimums
print min_76760_56840 >> minimums
print min_76760_59640 >> minimums
print min_76760_62440 >> minimums
print min_76760_65240 >> minimums
print min_76760_68040 >> minimums
print min_76760_70840 >> minimums
print min_76760_73640 >> minimums
print min_76760_76440 >> minimums
print min_76760_79240 >> minimums
print min_76760_82040 >> minimums
print min_76760_84840 >> minimums
print min_76760_87640 >> minimums
print min_77140_40040 >> minimums
print min_77140_42840 >> minimums
print min_77140_45640 >> minimums
print min_77140_48440 >> minimums
print min_77140_51240 >> minimums
print min_77140_54040 >> minimums
print min_77140_56840 >> minimums
print min_77140_59640 >> minimums
print min_77140_62440 >> minimums
print min_77140_65240 >> minimums
print min_77140_68040 >> minimums
print min_77140_70840 >> minimums
print min_77140_73640 >> minimums
print min_77140_76440 >> minimums
print min_77140_79240 >> minimums
print min_77140_82040 >> minimums
print min_77140_84840 >> minimums
print min_77140_87640 >> minimums
print min_77520_40040 >> minimums
print min_77520_42840 >> minimums
print min_77520_45640 >> minimums
print min_77520_48440 >> minimums
print min_77520_51240 >> minimums
print min_77520_54040 >> minimums
print min_77520_56840 >> minimums
print min_77520_59640 >> minimums
print min_77520_62440 >> minimums
print min_77520_65240 >> minimums
print min_77520_68040 >> minimums
print min_77520_70840 >> minimums
print min_77520_73640 >> minimums
print min_77520_76440 >> minimums
print min_77520_79240 >> minimums
print min_77520_82040 >> minimums
print min_77520_84840 >> minimums
print min_77520_87640 >> minimums
print min_77900_40040 >> minimums
print min_77900_42840 >> minimums
print min_77900_45640 >> minimums
print min_77900_48440 >> minimums
print min_77900_51240 >> minimums
print min_77900_54040 >> minimums
print min_77900_56840 >> minimums
print min_77900_59640 >> minimums
print min_77900_62440 >> minimums
print min_77900_65240 >> minimums
print min_77900_68040 >> minimums
print min_77900_70840 >> minimums
print min_77900_73640 >> minimums
print min_77900_76440 >> minimums
print min_77900_79240 >> minimums
print min_77900_82040 >> minimums
print min_77900_84840 >> minimums
print min_77900_87640 >> minimums
print min_78280_40040 >> minimums
print min_78280_42840 >> minimums
print min_78280_45640 >> minimums
print min_78280_48440 >> minimums
print min_78280_51240 >> minimums
print min_78280_54040 >> minimums
print min_78280_56840 >> minimums
print min_78280_59640 >> minimums
print min_78280_62440 >> minimums
print min_78280_65240 >> minimums
print min_78280_68040 >> minimums
print min_78280_70840 >> minimums
print min_78280_73640 >> minimums
print min_78280_76440 >> minimums
print min_78280_79240 >> minimums
print min_78280_82040 >> minimums
print min_78280_84840 >> minimums
print min_78280_87640 >> minimums
print min_78660_40040 >> minimums
print min_78660_42840 >> minimums
print min_78660_45640 >> minimums
print min_78660_48440 >> minimums
print min_78660_51240 >> minimums
print min_78660_54040 >> minimums
print min_78660_56840 >> minimums
print min_78660_59640 >> minimums
print min_78660_62440 >> minimums
print min_78660_65240 >> minimums
print min_78660_68040 >> minimums
print min_78660_70840 >> minimums
print min_78660_73640 >> minimums
print min_78660_76440 >> minimums
print min_78660_79240 >> minimums
print min_78660_82040 >> minimums
print min_78660_84840 >> minimums
print min_78660_87640 >> minimums
print min_79040_40040 >> minimums
print min_79040_42840 >> minimums
print min_79040_45640 >> minimums
print min_79040_48440 >> minimums
print min_79040_51240 >> minimums
print min_79040_54040 >> minimums
print min_79040_56840 >> minimums
print min_79040_59640 >> minimums
print min_79040_62440 >> minimums
print min_79040_65240 >> minimums
print min_79040_68040 >> minimums
print min_79040_70840 >> minimums
print min_79040_73640 >> minimums
print min_79040_76440 >> minimums
print min_79040_79240 >> minimums
print min_79040_82040 >> minimums
print min_79040_84840 >> minimums
print min_79040_87640 >> minimums
print min_80180_40040 >> minimums
print min_80180_42840 >> minimums
print min_80180_45640 >> minimums
print min_80180_48440 >> minimums
print min_80180_51240 >> minimums
print min_80180_54040 >> minimums
print min_80180_56840 >> minimums
print min_80180_59640 >> minimums
print min_80180_62440 >> minimums
print min_80180_65240 >> minimums
print min_80180_68040 >> minimums
print min_80180_70840 >> minimums
print min_80180_73640 >> minimums
print min_80180_76440 >> minimums
print min_80180_79240 >> minimums
print min_80180_82040 >> minimums
print min_80180_84840 >> minimums
print min_80180_87640 >> minimums
print min_80560_40040 >> minimums
print min_80560_42840 >> minimums
print min_80560_45640 >> minimums
print min_80560_48440 >> minimums
print min_80560_51240 >> minimums
print min_80560_54040 >> minimums
print min_80560_56840 >> minimums
print min_80560_59640 >> minimums
print min_80560_62440 >> minimums
print min_80560_65240 >> minimums
print min_80560_68040 >> minimums
print min_80560_70840 >> minimums
print min_80560_73640 >> minimums
print min_80560_76440 >> minimums
print min_80560_79240 >> minimums
print min_80560_82040 >> minimums
print min_80560_84840 >> minimums
print min_80560_87640 >> minimums
print min_80940_40040 >> minimums
print min_80940_42840 >> minimums
print min_80940_45640 >> minimums
print min_80940_48440 >> minimums
print min_80940_51240 >> minimums
print min_80940_54040 >> minimums
print min_80940_56840 >> minimums
print min_80940_59640 >> minimums
print min_80940_62440 >> minimums
print min_80940_65240 >> minimums
print min_80940_68040 >> minimums
print min_80940_70840 >> minimums
print min_80940_73640 >> minimums
print min_80940_76440 >> minimums
print min_80940_79240 >> minimums
print min_80940_82040 >> minimums
print min_80940_84840 >> minimums
print min_80940_87640 >> minimums
print min_81700_40040 >> minimums
print min_81700_42840 >> minimums
print min_81700_45640 >> minimums
print min_81700_48440 >> minimums
print min_81700_51240 >> minimums
print min_81700_54040 >> minimums
print min_81700_56840 >> minimums
print min_81700_59640 >> minimums
print min_81700_62440 >> minimums
print min_81700_65240 >> minimums
print min_81700_68040 >> minimums
print min_81700_70840 >> minimums
print min_81700_73640 >> minimums
print min_81700_76440 >> minimums
print min_81700_79240 >> minimums
print min_81700_82040 >> minimums
print min_81700_84840 >> minimums
print min_81700_87640 >> minimums
print min_82080_40040 >> minimums
print min_82080_42840 >> minimums
print min_82080_45640 >> minimums
print min_82080_48440 >> minimums
print min_82080_51240 >> minimums
print min_82080_54040 >> minimums
print min_82080_56840 >> minimums
print min_82080_59640 >> minimums
print min_82080_62440 >> minimums
print min_82080_65240 >> minimums
print min_82080_68040 >> minimums
print min_82080_70840 >> minimums
print min_82080_73640 >> minimums
print min_82080_76440 >> minimums
print min_82080_79240 >> minimums
print min_82080_82040 >> minimums
print min_82080_84840 >> minimums
print min_82080_87640 >> minimums
print min_83220_40040 >> minimums
print min_83220_42840 >> minimums
print min_83220_45640 >> minimums
print min_83220_48440 >> minimums
print min_83220_51240 >> minimums
print min_83220_54040 >> minimums
print min_83220_56840 >> minimums
print min_83220_59640 >> minimums
print min_83220_62440 >> minimums
print min_83220_65240 >> minimums
print min_83220_68040 >> minimums
print min_83220_70840 >> minimums
print min_83220_73640 >> minimums
print min_83220_76440 >> minimums
print min_83220_79240 >> minimums
print min_83220_82040 >> minimums
print min_83220_84840 >> minimums
print min_83220_87640 >> minimums
print min_83600_40040 >> minimums
print min_83600_42840 >> minimums
print min_83600_45640 >> minimums
print min_83600_48440 >> minimums
print min_83600_51240 >> minimums
print min_83600_54040 >> minimums
print min_83600_56840 >> minimums
print min_83600_59640 >> minimums
print min_83600_62440 >> minimums
print min_83600_65240 >> minimums
print min_83600_68040 >> minimums
print min_83600_70840 >> minimums
print min_83600_73640 >> minimums
print min_83600_76440 >> minimums
print min_83600_79240 >> minimums
print min_83600_82040 >> minimums
print min_83600_84840 >> minimums
print min_83600_87640 >> minimums
print min_84740_40040 >> minimums
print min_84740_42840 >> minimums
print min_84740_45640 >> minimums
print min_84740_48440 >> minimums
print min_84740_51240 >> minimums
print min_84740_54040 >> minimums
print min_84740_56840 >> minimums
print min_84740_59640 >> minimums
print min_84740_62440 >> minimums
print min_84740_65240 >> minimums
print min_84740_68040 >> minimums
print min_84740_70840 >> minimums
print min_84740_73640 >> minimums
print min_84740_76440 >> minimums
print min_84740_79240 >> minimums
print min_84740_82040 >> minimums
print min_84740_84840 >> minimums
print min_84740_87640 >> minimums
print min_85120_40040 >> minimums
print min_85120_42840 >> minimums
print min_85120_45640 >> minimums
print min_85120_48440 >> minimums
print min_85120_51240 >> minimums
print min_85120_54040 >> minimums
print min_85120_56840 >> minimums
print min_85120_59640 >> minimums
print min_85120_62440 >> minimums
print min_85120_65240 >> minimums
print min_85120_68040 >> minimums
print min_85120_70840 >> minimums
print min_85120_73640 >> minimums
print min_85120_76440 >> minimums
print min_85120_79240 >> minimums
print min_85120_82040 >> minimums
print min_85120_84840 >> minimums
print min_85120_87640 >> minimums
print min_85500_40040 >> minimums
print min_85500_42840 >> minimums
print min_85500_45640 >> minimums
print min_85500_48440 >> minimums
print min_85500_51240 >> minimums
print min_85500_54040 >> minimums
print min_85500_56840 >> minimums
print min_85500_59640 >> minimums
print min_85500_62440 >> minimums
print min_85500_65240 >> minimums
print min_85500_68040 >> minimums
print min_85500_70840 >> minimums
print min_85500_73640 >> minimums
print min_85500_76440 >> minimums
print min_85500_79240 >> minimums
print min_85500_82040 >> minimums
print min_85500_84840 >> minimums
print min_85500_87640 >> minimums
print min_85880_40040 >> minimums
print min_85880_42840 >> minimums
print min_85880_45640 >> minimums
print min_85880_48440 >> minimums
print min_85880_51240 >> minimums
print min_85880_54040 >> minimums
print min_85880_56840 >> minimums
print min_85880_59640 >> minimums
print min_85880_62440 >> minimums
print min_85880_65240 >> minimums
print min_85880_68040 >> minimums
print min_85880_70840 >> minimums
print min_85880_73640 >> minimums
print min_85880_76440 >> minimums
print min_85880_79240 >> minimums
print min_85880_82040 >> minimums
print min_85880_84840 >> minimums
print min_85880_87640 >> minimums
print min_86260_40040 >> minimums
print min_86260_42840 >> minimums
print min_86260_45640 >> minimums
print min_86260_48440 >> minimums
print min_86260_51240 >> minimums
print min_86260_54040 >> minimums
print min_86260_56840 >> minimums
print min_86260_59640 >> minimums
print min_86260_62440 >> minimums
print min_86260_65240 >> minimums
print min_86260_68040 >> minimums
print min_86260_70840 >> minimums
print min_86260_73640 >> minimums
print min_86260_76440 >> minimums
print min_86260_79240 >> minimums
print min_86260_82040 >> minimums
print min_86260_84840 >> minimums
print min_86260_87640 >> minimums
print min_87020_40040 >> minimums
print min_87020_42840 >> minimums
print min_87020_45640 >> minimums
print min_87020_48440 >> minimums
print min_87020_51240 >> minimums
print min_87020_54040 >> minimums
print min_87020_56840 >> minimums
print min_87020_59640 >> minimums
print min_87020_62440 >> minimums
print min_87020_65240 >> minimums
print min_87020_68040 >> minimums
print min_87020_70840 >> minimums
print min_87020_73640 >> minimums
print min_87020_76440 >> minimums
print min_87020_79240 >> minimums
print min_87020_82040 >> minimums
print min_87020_84840 >> minimums
print min_87020_87640 >> minimums
print min_87400_40040 >> minimums
print min_87400_42840 >> minimums
print min_87400_45640 >> minimums
print min_87400_48440 >> minimums
print min_87400_51240 >> minimums
print min_87400_54040 >> minimums
print min_87400_56840 >> minimums
print min_87400_59640 >> minimums
print min_87400_62440 >> minimums
print min_87400_65240 >> minimums
print min_87400_68040 >> minimums
print min_87400_70840 >> minimums
print min_87400_73640 >> minimums
print min_87400_76440 >> minimums
print min_87400_79240 >> minimums
print min_87400_82040 >> minimums
print min_87400_84840 >> minimums
print min_87400_87640 >> minimums
print min_87780_40040 >> minimums
print min_87780_42840 >> minimums
print min_87780_45640 >> minimums
print min_87780_48440 >> minimums
print min_87780_51240 >> minimums
print min_87780_54040 >> minimums
print min_87780_56840 >> minimums
print min_87780_59640 >> minimums
print min_87780_62440 >> minimums
print min_87780_65240 >> minimums
print min_87780_68040 >> minimums
print min_87780_70840 >> minimums
print min_87780_73640 >> minimums
print min_87780_76440 >> minimums
print min_87780_79240 >> minimums
print min_87780_82040 >> minimums
print min_87780_84840 >> minimums
print min_87780_87640 >> minimums
print min_88160_40040 >> minimums
print min_88160_42840 >> minimums
print min_88160_45640 >> minimums
print min_88160_48440 >> minimums
print min_88160_51240 >> minimums
print min_88160_54040 >> minimums
print min_88160_56840 >> minimums
print min_88160_59640 >> minimums
print min_88160_62440 >> minimums
print min_88160_65240 >> minimums
print min_88160_68040 >> minimums
print min_88160_70840 >> minimums
print min_88160_73640 >> minimums
print min_88160_76440 >> minimums
print min_88160_79240 >> minimums
print min_88160_82040 >> minimums
print min_88160_84840 >> minimums
print min_88160_87640 >> minimums
print min_88540_40040 >> minimums
print min_88540_42840 >> minimums
print min_88540_45640 >> minimums
print min_88540_48440 >> minimums
print min_88540_51240 >> minimums
print min_88540_54040 >> minimums
print min_88540_56840 >> minimums
print min_88540_59640 >> minimums
print min_88540_62440 >> minimums
print min_88540_65240 >> minimums
print min_88540_68040 >> minimums
print min_88540_70840 >> minimums
print min_88540_73640 >> minimums
print min_88540_76440 >> minimums
print min_88540_79240 >> minimums
print min_88540_82040 >> minimums
print min_88540_84840 >> minimums
print min_88540_87640 >> minimums
print min_88920_40040 >> minimums
print min_88920_42840 >> minimums
print min_88920_45640 >> minimums
print min_88920_48440 >> minimums
print min_88920_51240 >> minimums
print min_88920_54040 >> minimums
print min_88920_56840 >> minimums
print min_88920_59640 >> minimums
print min_88920_62440 >> minimums
print min_88920_65240 >> minimums
print min_88920_68040 >> minimums
print min_88920_70840 >> minimums
print min_88920_73640 >> minimums
print min_88920_76440 >> minimums
print min_88920_79240 >> minimums
print min_88920_82040 >> minimums
print min_88920_84840 >> minimums
print min_88920_87640 >> minimums
print min_89300_40040 >> minimums
print min_89300_42840 >> minimums
print min_89300_45640 >> minimums
print min_89300_48440 >> minimums
print min_89300_51240 >> minimums
print min_89300_54040 >> minimums
print min_89300_56840 >> minimums
print min_89300_59640 >> minimums
print min_89300_62440 >> minimums
print min_89300_65240 >> minimums
print min_89300_68040 >> minimums
print min_89300_70840 >> minimums
print min_89300_73640 >> minimums
print min_89300_76440 >> minimums
print min_89300_79240 >> minimums
print min_89300_82040 >> minimums
print min_89300_84840 >> minimums
print min_89300_87640 >> minimums
print min_90060_40040 >> minimums
print min_90060_42840 >> minimums
print min_90060_45640 >> minimums
print min_90060_48440 >> minimums
print min_90060_51240 >> minimums
print min_90060_54040 >> minimums
print min_90060_56840 >> minimums
print min_90060_59640 >> minimums
print min_90060_62440 >> minimums
print min_90060_65240 >> minimums
print min_90060_68040 >> minimums
print min_90060_70840 >> minimums
print min_90060_73640 >> minimums
print min_90060_76440 >> minimums
print min_90060_79240 >> minimums
print min_90060_82040 >> minimums
print min_90060_84840 >> minimums
print min_90060_87640 >> minimums
print min_90440_40040 >> minimums
print min_90440_42840 >> minimums
print min_90440_45640 >> minimums
print min_90440_48440 >> minimums
print min_90440_51240 >> minimums
print min_90440_54040 >> minimums
print min_90440_56840 >> minimums
print min_90440_59640 >> minimums
print min_90440_62440 >> minimums
print min_90440_65240 >> minimums
print min_90440_68040 >> minimums
print min_90440_70840 >> minimums
print min_90440_73640 >> minimums
print min_90440_76440 >> minimums
print min_90440_79240 >> minimums
print min_90440_82040 >> minimums
print min_90440_84840 >> minimums
print min_90440_87640 >> minimums
print min_90820_40040 >> minimums
print min_90820_42840 >> minimums
print min_90820_45640 >> minimums
print min_90820_48440 >> minimums
print min_90820_51240 >> minimums
print min_90820_54040 >> minimums
print min_90820_56840 >> minimums
print min_90820_59640 >> minimums
print min_90820_62440 >> minimums
print min_90820_65240 >> minimums
print min_90820_68040 >> minimums
print min_90820_70840 >> minimums
print min_90820_73640 >> minimums
print min_90820_76440 >> minimums
print min_90820_79240 >> minimums
print min_90820_82040 >> minimums
print min_90820_84840 >> minimums
print min_90820_87640 >> minimums
print min_91200_40040 >> minimums
print min_91200_42840 >> minimums
print min_91200_45640 >> minimums
print min_91200_48440 >> minimums
print min_91200_51240 >> minimums
print min_91200_54040 >> minimums
print min_91200_56840 >> minimums
print min_91200_59640 >> minimums
print min_91200_62440 >> minimums
print min_91200_65240 >> minimums
print min_91200_68040 >> minimums
print min_91200_70840 >> minimums
print min_91200_73640 >> minimums
print min_91200_76440 >> minimums
print min_91200_79240 >> minimums
print min_91200_82040 >> minimums
print min_91200_84840 >> minimums
print min_91200_87640 >> minimums
print min_91580_40040 >> minimums
print min_91580_42840 >> minimums
print min_91580_45640 >> minimums
print min_91580_48440 >> minimums
print min_91580_51240 >> minimums
print min_91580_54040 >> minimums
print min_91580_56840 >> minimums
print min_91580_59640 >> minimums
print min_91580_62440 >> minimums
print min_91580_65240 >> minimums
print min_91580_68040 >> minimums
print min_91580_70840 >> minimums
print min_91580_73640 >> minimums
print min_91580_76440 >> minimums
print min_91580_79240 >> minimums
print min_91580_82040 >> minimums
print min_91580_84840 >> minimums
print min_91580_87640 >> minimums
print min_91960_40040 >> minimums
print min_91960_42840 >> minimums
print min_91960_45640 >> minimums
print min_91960_48440 >> minimums
print min_91960_51240 >> minimums
print min_91960_54040 >> minimums
print min_91960_56840 >> minimums
print min_91960_59640 >> minimums
print min_91960_62440 >> minimums
print min_91960_65240 >> minimums
print min_91960_68040 >> minimums
print min_91960_70840 >> minimums
print min_91960_73640 >> minimums
print min_91960_76440 >> minimums
print min_91960_79240 >> minimums
print min_91960_82040 >> minimums
print min_91960_84840 >> minimums
print min_91960_87640 >> minimums
print min_92340_40040 >> minimums
print min_92340_42840 >> minimums
print min_92340_45640 >> minimums
print min_92340_48440 >> minimums
print min_92340_51240 >> minimums
print min_92340_54040 >> minimums
print min_92340_56840 >> minimums
print min_92340_59640 >> minimums
print min_92340_62440 >> minimums
print min_92340_65240 >> minimums
print min_92340_68040 >> minimums
print min_92340_70840 >> minimums
print min_92340_73640 >> minimums
print min_92340_76440 >> minimums
print min_92340_79240 >> minimums
print min_92340_82040 >> minimums
print min_92340_84840 >> minimums
print min_92340_87640 >> minimums
print min_92720_40040 >> minimums
print min_92720_42840 >> minimums
print min_92720_45640 >> minimums
print min_92720_48440 >> minimums
print min_92720_51240 >> minimums
print min_92720_54040 >> minimums
print min_92720_56840 >> minimums
print min_92720_59640 >> minimums
print min_92720_62440 >> minimums
print min_92720_65240 >> minimums
print min_92720_68040 >> minimums
print min_92720_70840 >> minimums
print min_92720_73640 >> minimums
print min_92720_76440 >> minimums
print min_92720_79240 >> minimums
print min_92720_82040 >> minimums
print min_92720_84840 >> minimums
print min_92720_87640 >> minimums
print min_93100_40040 >> minimums
print min_93100_42840 >> minimums
print min_93100_45640 >> minimums
print min_93100_48440 >> minimums
print min_93100_51240 >> minimums
print min_93100_54040 >> minimums
print min_93100_56840 >> minimums
print min_93100_59640 >> minimums
print min_93100_62440 >> minimums
print min_93100_65240 >> minimums
print min_93100_68040 >> minimums
print min_93100_70840 >> minimums
print min_93100_73640 >> minimums
print min_93100_76440 >> minimums
print min_93100_79240 >> minimums
print min_93100_82040 >> minimums
print min_93100_84840 >> minimums
print min_93100_87640 >> minimums
print min_93480_40040 >> minimums
print min_93480_42840 >> minimums
print min_93480_45640 >> minimums
print min_93480_48440 >> minimums
print min_93480_51240 >> minimums
print min_93480_54040 >> minimums
print min_93480_56840 >> minimums
print min_93480_59640 >> minimums
print min_93480_62440 >> minimums
print min_93480_65240 >> minimums
print min_93480_68040 >> minimums
print min_93480_70840 >> minimums
print min_93480_73640 >> minimums
print min_93480_76440 >> minimums
print min_93480_79240 >> minimums
print min_93480_82040 >> minimums
print min_93480_84840 >> minimums
print min_93480_87640 >> minimums

exit
.endc