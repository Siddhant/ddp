.title 1-layer Power Grid for b01.points
* resistance segment model:
.subckt Rseg 1 3
R1 1 2 0.583
L1 2 3 0.003n
C1 1 0 0.25e-12
C2 3 0 0.25e-12
.ends
* the horizontal resistors:
X1 n_40660_40040 n_41040_40040 Rseg
X2 n_41040_40040 n_42180_40040 Rseg
X3 n_42180_40040 n_42560_40040 Rseg
X4 n_42560_40040 n_42940_40040 Rseg
X5 n_42940_40040 n_43700_40040 Rseg
X6 n_43700_40040 n_44080_40040 Rseg
X7 n_44080_40040 n_44840_40040 Rseg
X8 n_44840_40040 n_45220_40040 Rseg
X9 n_45220_40040 n_45600_40040 Rseg
X10 n_45600_40040 n_46360_40040 Rseg
X11 n_46360_40040 n_46740_40040 Rseg
X12 n_46740_40040 n_47120_40040 Rseg
X13 n_47120_40040 n_47500_40040 Rseg
X14 n_47500_40040 n_47880_40040 Rseg
X15 n_47880_40040 n_48260_40040 Rseg
X16 n_48260_40040 n_48640_40040 Rseg
X17 n_48640_40040 n_49400_40040 Rseg
X18 n_49400_40040 n_49780_40040 Rseg
X19 n_49780_40040 n_50160_40040 Rseg
X20 n_50160_40040 n_50540_40040 Rseg
X21 n_50540_40040 n_51300_40040 Rseg
X22 n_51300_40040 n_51680_40040 Rseg
X23 n_51680_40040 n_52440_40040 Rseg
X24 n_52440_40040 n_52820_40040 Rseg
X25 n_52820_40040 n_53580_40040 Rseg
X26 n_53580_40040 n_53960_40040 Rseg
X27 n_53960_40040 n_54340_40040 Rseg
X28 n_54340_40040 n_54720_40040 Rseg
X29 n_54720_40040 n_55100_40040 Rseg
X30 n_40660_42840 n_41040_42840 Rseg
X31 n_41040_42840 n_42180_42840 Rseg
X32 n_42180_42840 n_42560_42840 Rseg
X33 n_42560_42840 n_42940_42840 Rseg
X34 n_42940_42840 n_43700_42840 Rseg
X35 n_43700_42840 n_44080_42840 Rseg
X36 n_44080_42840 n_44840_42840 Rseg
X37 n_44840_42840 n_45220_42840 Rseg
X38 n_45220_42840 n_45600_42840 Rseg
X39 n_45600_42840 n_46360_42840 Rseg
X40 n_46360_42840 n_46740_42840 Rseg
X41 n_46740_42840 n_47120_42840 Rseg
X42 n_47120_42840 n_47500_42840 Rseg
X43 n_47500_42840 n_47880_42840 Rseg
X44 n_47880_42840 n_48260_42840 Rseg
X45 n_48260_42840 n_48640_42840 Rseg
X46 n_48640_42840 n_49400_42840 Rseg
X47 n_49400_42840 n_49780_42840 Rseg
X48 n_49780_42840 n_50160_42840 Rseg
X49 n_50160_42840 n_50540_42840 Rseg
X50 n_50540_42840 n_51300_42840 Rseg
X51 n_51300_42840 n_51680_42840 Rseg
X52 n_51680_42840 n_52440_42840 Rseg
X53 n_52440_42840 n_52820_42840 Rseg
X54 n_52820_42840 n_53580_42840 Rseg
X55 n_53580_42840 n_53960_42840 Rseg
X56 n_53960_42840 n_54340_42840 Rseg
X57 n_54340_42840 n_54720_42840 Rseg
X58 n_54720_42840 n_55100_42840 Rseg
X59 n_40660_45640 n_41040_45640 Rseg
X60 n_41040_45640 n_42180_45640 Rseg
X61 n_42180_45640 n_42560_45640 Rseg
X62 n_42560_45640 n_42940_45640 Rseg
X63 n_42940_45640 n_43700_45640 Rseg
X64 n_43700_45640 n_44080_45640 Rseg
X65 n_44080_45640 n_44840_45640 Rseg
X66 n_44840_45640 n_45220_45640 Rseg
X67 n_45220_45640 n_45600_45640 Rseg
X68 n_45600_45640 n_46360_45640 Rseg
X69 n_46360_45640 n_46740_45640 Rseg
X70 n_46740_45640 n_47120_45640 Rseg
X71 n_47120_45640 n_47500_45640 Rseg
X72 n_47500_45640 n_47880_45640 Rseg
X73 n_47880_45640 n_48260_45640 Rseg
X74 n_48260_45640 n_48640_45640 Rseg
X75 n_48640_45640 n_49400_45640 Rseg
X76 n_49400_45640 n_49780_45640 Rseg
X77 n_49780_45640 n_50160_45640 Rseg
X78 n_50160_45640 n_50540_45640 Rseg
X79 n_50540_45640 n_51300_45640 Rseg
X80 n_51300_45640 n_51680_45640 Rseg
X81 n_51680_45640 n_52440_45640 Rseg
X82 n_52440_45640 n_52820_45640 Rseg
X83 n_52820_45640 n_53580_45640 Rseg
X84 n_53580_45640 n_53960_45640 Rseg
X85 n_53960_45640 n_54340_45640 Rseg
X86 n_54340_45640 n_54720_45640 Rseg
X87 n_54720_45640 n_55100_45640 Rseg
X88 n_40660_48440 n_41040_48440 Rseg
X89 n_41040_48440 n_42180_48440 Rseg
X90 n_42180_48440 n_42560_48440 Rseg
X91 n_42560_48440 n_42940_48440 Rseg
X92 n_42940_48440 n_43700_48440 Rseg
X93 n_43700_48440 n_44080_48440 Rseg
X94 n_44080_48440 n_44840_48440 Rseg
X95 n_44840_48440 n_45220_48440 Rseg
X96 n_45220_48440 n_45600_48440 Rseg
X97 n_45600_48440 n_46360_48440 Rseg
X98 n_46360_48440 n_46740_48440 Rseg
X99 n_46740_48440 n_47120_48440 Rseg
X100 n_47120_48440 n_47500_48440 Rseg
X101 n_47500_48440 n_47880_48440 Rseg
X102 n_47880_48440 n_48260_48440 Rseg
X103 n_48260_48440 n_48640_48440 Rseg
X104 n_48640_48440 n_49400_48440 Rseg
X105 n_49400_48440 n_49780_48440 Rseg
X106 n_49780_48440 n_50160_48440 Rseg
X107 n_50160_48440 n_50540_48440 Rseg
X108 n_50540_48440 n_51300_48440 Rseg
X109 n_51300_48440 n_51680_48440 Rseg
X110 n_51680_48440 n_52440_48440 Rseg
X111 n_52440_48440 n_52820_48440 Rseg
X112 n_52820_48440 n_53580_48440 Rseg
X113 n_53580_48440 n_53960_48440 Rseg
X114 n_53960_48440 n_54340_48440 Rseg
X115 n_54340_48440 n_54720_48440 Rseg
X116 n_54720_48440 n_55100_48440 Rseg
X117 n_40660_51240 n_41040_51240 Rseg
X118 n_41040_51240 n_42180_51240 Rseg
X119 n_42180_51240 n_42560_51240 Rseg
X120 n_42560_51240 n_42940_51240 Rseg
X121 n_42940_51240 n_43700_51240 Rseg
X122 n_43700_51240 n_44080_51240 Rseg
X123 n_44080_51240 n_44840_51240 Rseg
X124 n_44840_51240 n_45220_51240 Rseg
X125 n_45220_51240 n_45600_51240 Rseg
X126 n_45600_51240 n_46360_51240 Rseg
X127 n_46360_51240 n_46740_51240 Rseg
X128 n_46740_51240 n_47120_51240 Rseg
X129 n_47120_51240 n_47500_51240 Rseg
X130 n_47500_51240 n_47880_51240 Rseg
X131 n_47880_51240 n_48260_51240 Rseg
X132 n_48260_51240 n_48640_51240 Rseg
X133 n_48640_51240 n_49400_51240 Rseg
X134 n_49400_51240 n_49780_51240 Rseg
X135 n_49780_51240 n_50160_51240 Rseg
X136 n_50160_51240 n_50540_51240 Rseg
X137 n_50540_51240 n_51300_51240 Rseg
X138 n_51300_51240 n_51680_51240 Rseg
X139 n_51680_51240 n_52440_51240 Rseg
X140 n_52440_51240 n_52820_51240 Rseg
X141 n_52820_51240 n_53580_51240 Rseg
X142 n_53580_51240 n_53960_51240 Rseg
X143 n_53960_51240 n_54340_51240 Rseg
X144 n_54340_51240 n_54720_51240 Rseg
X145 n_54720_51240 n_55100_51240 Rseg
* the vertical resistors:
X146 n_40660_40040 n_40660_42840 Rseg
X147 n_40660_42840 n_40660_45640 Rseg
X148 n_40660_45640 n_40660_48440 Rseg
X149 n_40660_48440 n_40660_51240 Rseg
X150 n_41040_40040 n_41040_42840 Rseg
X151 n_41040_42840 n_41040_45640 Rseg
X152 n_41040_45640 n_41040_48440 Rseg
X153 n_41040_48440 n_41040_51240 Rseg
X154 n_42180_40040 n_42180_42840 Rseg
X155 n_42180_42840 n_42180_45640 Rseg
X156 n_42180_45640 n_42180_48440 Rseg
X157 n_42180_48440 n_42180_51240 Rseg
X158 n_42560_40040 n_42560_42840 Rseg
X159 n_42560_42840 n_42560_45640 Rseg
X160 n_42560_45640 n_42560_48440 Rseg
X161 n_42560_48440 n_42560_51240 Rseg
X162 n_42940_40040 n_42940_42840 Rseg
X163 n_42940_42840 n_42940_45640 Rseg
X164 n_42940_45640 n_42940_48440 Rseg
X165 n_42940_48440 n_42940_51240 Rseg
X166 n_43700_40040 n_43700_42840 Rseg
X167 n_43700_42840 n_43700_45640 Rseg
X168 n_43700_45640 n_43700_48440 Rseg
X169 n_43700_48440 n_43700_51240 Rseg
X170 n_44080_40040 n_44080_42840 Rseg
X171 n_44080_42840 n_44080_45640 Rseg
X172 n_44080_45640 n_44080_48440 Rseg
X173 n_44080_48440 n_44080_51240 Rseg
X174 n_44840_40040 n_44840_42840 Rseg
X175 n_44840_42840 n_44840_45640 Rseg
X176 n_44840_45640 n_44840_48440 Rseg
X177 n_44840_48440 n_44840_51240 Rseg
X178 n_45220_40040 n_45220_42840 Rseg
X179 n_45220_42840 n_45220_45640 Rseg
X180 n_45220_45640 n_45220_48440 Rseg
X181 n_45220_48440 n_45220_51240 Rseg
X182 n_45600_40040 n_45600_42840 Rseg
X183 n_45600_42840 n_45600_45640 Rseg
X184 n_45600_45640 n_45600_48440 Rseg
X185 n_45600_48440 n_45600_51240 Rseg
X186 n_46360_40040 n_46360_42840 Rseg
X187 n_46360_42840 n_46360_45640 Rseg
X188 n_46360_45640 n_46360_48440 Rseg
X189 n_46360_48440 n_46360_51240 Rseg
X190 n_46740_40040 n_46740_42840 Rseg
X191 n_46740_42840 n_46740_45640 Rseg
X192 n_46740_45640 n_46740_48440 Rseg
X193 n_46740_48440 n_46740_51240 Rseg
X194 n_47120_40040 n_47120_42840 Rseg
X195 n_47120_42840 n_47120_45640 Rseg
X196 n_47120_45640 n_47120_48440 Rseg
X197 n_47120_48440 n_47120_51240 Rseg
X198 n_47500_40040 n_47500_42840 Rseg
X199 n_47500_42840 n_47500_45640 Rseg
X200 n_47500_45640 n_47500_48440 Rseg
X201 n_47500_48440 n_47500_51240 Rseg
X202 n_47880_40040 n_47880_42840 Rseg
X203 n_47880_42840 n_47880_45640 Rseg
X204 n_47880_45640 n_47880_48440 Rseg
X205 n_47880_48440 n_47880_51240 Rseg
X206 n_48260_40040 n_48260_42840 Rseg
X207 n_48260_42840 n_48260_45640 Rseg
X208 n_48260_45640 n_48260_48440 Rseg
X209 n_48260_48440 n_48260_51240 Rseg
X210 n_48640_40040 n_48640_42840 Rseg
X211 n_48640_42840 n_48640_45640 Rseg
X212 n_48640_45640 n_48640_48440 Rseg
X213 n_48640_48440 n_48640_51240 Rseg
X214 n_49400_40040 n_49400_42840 Rseg
X215 n_49400_42840 n_49400_45640 Rseg
X216 n_49400_45640 n_49400_48440 Rseg
X217 n_49400_48440 n_49400_51240 Rseg
X218 n_49780_40040 n_49780_42840 Rseg
X219 n_49780_42840 n_49780_45640 Rseg
X220 n_49780_45640 n_49780_48440 Rseg
X221 n_49780_48440 n_49780_51240 Rseg
X222 n_50160_40040 n_50160_42840 Rseg
X223 n_50160_42840 n_50160_45640 Rseg
X224 n_50160_45640 n_50160_48440 Rseg
X225 n_50160_48440 n_50160_51240 Rseg
X226 n_50540_40040 n_50540_42840 Rseg
X227 n_50540_42840 n_50540_45640 Rseg
X228 n_50540_45640 n_50540_48440 Rseg
X229 n_50540_48440 n_50540_51240 Rseg
X230 n_51300_40040 n_51300_42840 Rseg
X231 n_51300_42840 n_51300_45640 Rseg
X232 n_51300_45640 n_51300_48440 Rseg
X233 n_51300_48440 n_51300_51240 Rseg
X234 n_51680_40040 n_51680_42840 Rseg
X235 n_51680_42840 n_51680_45640 Rseg
X236 n_51680_45640 n_51680_48440 Rseg
X237 n_51680_48440 n_51680_51240 Rseg
X238 n_52440_40040 n_52440_42840 Rseg
X239 n_52440_42840 n_52440_45640 Rseg
X240 n_52440_45640 n_52440_48440 Rseg
X241 n_52440_48440 n_52440_51240 Rseg
X242 n_52820_40040 n_52820_42840 Rseg
X243 n_52820_42840 n_52820_45640 Rseg
X244 n_52820_45640 n_52820_48440 Rseg
X245 n_52820_48440 n_52820_51240 Rseg
X246 n_53580_40040 n_53580_42840 Rseg
X247 n_53580_42840 n_53580_45640 Rseg
X248 n_53580_45640 n_53580_48440 Rseg
X249 n_53580_48440 n_53580_51240 Rseg
X250 n_53960_40040 n_53960_42840 Rseg
X251 n_53960_42840 n_53960_45640 Rseg
X252 n_53960_45640 n_53960_48440 Rseg
X253 n_53960_48440 n_53960_51240 Rseg
X254 n_54340_40040 n_54340_42840 Rseg
X255 n_54340_42840 n_54340_45640 Rseg
X256 n_54340_45640 n_54340_48440 Rseg
X257 n_54340_48440 n_54340_51240 Rseg
X258 n_54720_40040 n_54720_42840 Rseg
X259 n_54720_42840 n_54720_45640 Rseg
X260 n_54720_45640 n_54720_48440 Rseg
X261 n_54720_48440 n_54720_51240 Rseg
X262 n_55100_40040 n_55100_42840 Rseg
X263 n_55100_42840 n_55100_45640 Rseg
X264 n_55100_45640 n_55100_48440 Rseg
X265 n_55100_48440 n_55100_51240 Rseg
* voltage source is placed at (x_min, y_min)
Vin n_40660_40040 0 DC 1.0

I1 n_40660_48440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I2 n_55100_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I3 n_40660_51240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I4 n_42180_51240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I5 n_44080_48440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I6 n_45220_48440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I7 n_50540_48440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I8 n_41040_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I9 n_53960_48440 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I10 n_52440_51240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I11 n_45600_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I12 n_44080_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I13 n_44080_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I14 n_42180_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I15 n_44080_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I16 n_42940_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I17 n_47500_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I18 n_53960_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I19 n_54720_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I20 n_51300_51240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I21 n_50160_51240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I22 n_43700_51240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I23 n_47880_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I24 n_54340_51240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I25 n_53580_51240 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I26 n_55100_51240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I27 n_51300_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I28 n_55100_48440 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I29 n_48260_45640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I30 n_48260_51240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I31 n_50540_42840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I32 n_45600_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I33 n_44080_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I34 n_42560_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I35 n_40660_42840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I36 n_47120_42840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I37 n_49780_42840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I38 n_49400_45640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I39 n_50540_45640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I40 n_54720_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I41 n_54720_45640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I42 n_51300_51240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I43 n_50160_51240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I44 n_49400_51240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I45 n_43700_51240 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I46 n_52440_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I47 n_46740_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I48 n_40660_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I49 n_48260_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I50 n_40660_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I51 n_42180_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I52 n_44080_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I53 n_45220_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I54 n_41040_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I55 n_48260_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I56 n_53960_48440 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I57 n_52440_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I58 n_48260_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I59 n_50160_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I60 n_45600_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I61 n_44080_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I62 n_42560_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I63 n_42180_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I64 n_40660_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I65 n_44080_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I66 n_42940_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I67 n_47500_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I68 n_54720_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I69 n_54720_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I70 n_51300_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I71 n_50160_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I72 n_49400_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I73 n_43700_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I74 n_52440_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I75 n_46740_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I76 n_47880_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I77 n_53580_51240 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I78 n_55100_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I79 n_42180_48440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I80 n_42180_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I81 n_44840_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I82 n_41040_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I83 n_53960_48440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I84 n_52440_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I85 n_48260_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I86 n_42180_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I87 n_44080_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I88 n_42940_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I89 n_53960_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I90 n_54720_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I91 n_51300_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I92 n_50160_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I93 n_49400_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I94 n_43700_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I95 n_46360_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I96 n_46740_48440 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I97 n_47880_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I98 n_53580_51240 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I99 n_40660_48440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I100 n_48260_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I101 n_55100_42840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I102 n_55100_51240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I103 n_51300_48440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I104 n_55100_48440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I105 n_40660_51240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I106 n_42180_48440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I107 n_44840_45640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I108 n_44080_48440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I109 n_45220_48440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I110 n_48260_51240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I111 n_50160_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I112 n_50540_42840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I113 n_47120_42840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I114 n_49780_42840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I115 n_49400_45640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I116 n_50540_45640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I117 n_47500_45640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I118 n_53960_42840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I119 n_54720_45640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I120 n_51300_51240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I121 n_50160_51240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I122 n_49400_51240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I123 n_43700_51240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I124 n_46360_51240 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I125 n_46740_48440 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I126 n_40660_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I127 n_48260_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I128 n_55100_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I129 n_51300_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I130 n_55100_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I131 n_40660_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I132 n_42180_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I133 n_44840_45640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I134 n_44080_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I135 n_45220_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I136 n_48260_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I137 n_50160_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I138 n_50540_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I139 n_47500_45640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I140 n_47120_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I141 n_50160_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I142 n_49400_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I143 n_46360_51240 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I144 n_46740_48440 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I145 n_40660_48440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I146 n_48260_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I147 n_55100_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I148 n_55100_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I149 n_51300_48440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I150 n_55100_48440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I151 n_40660_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I152 n_42180_48440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I153 n_41040_45640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I154 n_53960_48440 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I155 n_52440_45640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I156 n_50160_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I157 n_45600_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I158 n_44080_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I159 n_44080_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I160 n_44080_45640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I161 n_42940_45640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I162 n_53960_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I163 n_54720_45640 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I164 n_51300_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I165 n_47120_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I166 n_43700_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I167 n_47880_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I168 n_54340_51240 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I169 n_48260_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I170 n_55100_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I171 n_50160_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I172 n_45600_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I173 n_44080_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I174 n_44080_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I175 n_47120_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I176 n_49780_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I177 n_49400_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I178 n_50540_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I179 n_53960_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I180 n_54720_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I181 n_51300_51240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I182 n_47120_51240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I183 n_43700_51240 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I184 n_40660_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I185 n_40660_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I186 n_42180_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I187 n_44840_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I188 n_41040_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I189 n_53960_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I190 n_52440_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I191 n_48260_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I192 n_44080_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I193 n_42940_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I194 n_47120_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I195 n_50160_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I196 n_49400_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I197 n_43700_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I198 n_46360_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I199 n_46740_48440 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I200 n_47880_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I201 n_54340_51240 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I202 n_40660_48440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I203 n_55100_42840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I204 n_55100_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I205 n_51300_48440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I206 n_55100_48440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I207 n_40660_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I208 n_42180_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I209 n_44080_48440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I210 n_45220_48440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I211 n_47880_48440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I212 n_50540_48440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I213 n_48260_45640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I214 n_53960_48440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I215 n_48260_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I216 n_52440_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I217 n_42180_42840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I218 n_40660_42840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I219 n_49400_48440 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I220 n_50540_45640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I221 n_47500_45640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I222 n_53960_42840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I223 n_54720_45640 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I224 n_51300_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I225 n_50160_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I226 n_49400_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I227 n_43700_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I228 n_47880_42840 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I229 n_54340_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I230 n_53580_51240 0 PWL(18000ps 0uA 18030ps 0uA 18031ps 30uA 18059ps 30uA 18060ps 0uA)
I231 n_52820_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I232 n_55100_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I233 n_45600_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I234 n_44840_45640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I235 n_47880_48440 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I236 n_41040_45640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I237 n_48260_45640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I238 n_42180_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I239 n_40660_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I240 n_47120_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I241 n_53960_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I242 n_54720_40040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I243 n_43700_51240 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I244 n_52440_40040 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I245 n_51680_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I246 n_48640_42840 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I247 n_45600_45640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I248 n_46360_45640 0 PWL(20000ps 0uA 20030ps 0uA 20031ps 30uA 20059ps 30uA 20060ps 0uA)
I249 n_52820_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I250 n_40660_48440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I251 n_48260_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I252 n_55100_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I253 n_55100_51240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I254 n_45600_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I255 n_51300_48440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I256 n_55100_48440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I257 n_40660_51240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I258 n_42180_48440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I259 n_50540_48440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I260 n_41040_45640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I261 n_48260_45640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I262 n_52440_45640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I263 n_52440_51240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I264 n_50160_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I265 n_45600_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I266 n_44080_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I267 n_42560_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I268 n_40660_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I269 n_47120_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I270 n_49400_48440 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I271 n_50540_45640 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I272 n_53960_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I273 n_54720_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I274 n_43700_51240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I275 n_52440_40040 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I276 n_51680_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I277 n_48640_42840 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I278 n_53580_51240 0 PWL(22000ps 0uA 22030ps 0uA 22031ps 30uA 22059ps 30uA 22060ps 0uA)
I279 n_40660_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I280 n_40660_51240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I281 n_42180_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I282 n_44840_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I283 n_47880_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I284 n_50540_48440 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I285 n_41040_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I286 n_48260_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I287 n_52440_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I288 n_48260_51240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I289 n_52440_51240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I290 n_50540_42840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I291 n_45600_40040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I292 n_44080_40040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I293 n_42560_40040 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I294 n_42180_42840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I295 n_40660_42840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I296 n_44080_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I297 n_42940_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I298 n_49780_42840 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I299 n_49400_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I300 n_50540_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I301 n_47500_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I302 n_49400_51240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I303 n_53580_51240 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I304 n_45600_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
I305 n_46360_45640 0 PWL(24000ps 0uA 24030ps 0uA 24031ps 30uA 24059ps 30uA 24060ps 0uA)
.tran 1ps 28000ps
.control
run
* calculate minimum value of voltage at each node:
let min_40660_40040 = minimum(v(n_40660_40040))
let min_40660_42840 = minimum(v(n_40660_42840))
let min_40660_45640 = minimum(v(n_40660_45640))
let min_40660_48440 = minimum(v(n_40660_48440))
let min_40660_51240 = minimum(v(n_40660_51240))
let min_41040_40040 = minimum(v(n_41040_40040))
let min_41040_42840 = minimum(v(n_41040_42840))
let min_41040_45640 = minimum(v(n_41040_45640))
let min_41040_48440 = minimum(v(n_41040_48440))
let min_41040_51240 = minimum(v(n_41040_51240))
let min_42180_40040 = minimum(v(n_42180_40040))
let min_42180_42840 = minimum(v(n_42180_42840))
let min_42180_45640 = minimum(v(n_42180_45640))
let min_42180_48440 = minimum(v(n_42180_48440))
let min_42180_51240 = minimum(v(n_42180_51240))
let min_42560_40040 = minimum(v(n_42560_40040))
let min_42560_42840 = minimum(v(n_42560_42840))
let min_42560_45640 = minimum(v(n_42560_45640))
let min_42560_48440 = minimum(v(n_42560_48440))
let min_42560_51240 = minimum(v(n_42560_51240))
let min_42940_40040 = minimum(v(n_42940_40040))
let min_42940_42840 = minimum(v(n_42940_42840))
let min_42940_45640 = minimum(v(n_42940_45640))
let min_42940_48440 = minimum(v(n_42940_48440))
let min_42940_51240 = minimum(v(n_42940_51240))
let min_43700_40040 = minimum(v(n_43700_40040))
let min_43700_42840 = minimum(v(n_43700_42840))
let min_43700_45640 = minimum(v(n_43700_45640))
let min_43700_48440 = minimum(v(n_43700_48440))
let min_43700_51240 = minimum(v(n_43700_51240))
let min_44080_40040 = minimum(v(n_44080_40040))
let min_44080_42840 = minimum(v(n_44080_42840))
let min_44080_45640 = minimum(v(n_44080_45640))
let min_44080_48440 = minimum(v(n_44080_48440))
let min_44080_51240 = minimum(v(n_44080_51240))
let min_44840_40040 = minimum(v(n_44840_40040))
let min_44840_42840 = minimum(v(n_44840_42840))
let min_44840_45640 = minimum(v(n_44840_45640))
let min_44840_48440 = minimum(v(n_44840_48440))
let min_44840_51240 = minimum(v(n_44840_51240))
let min_45220_40040 = minimum(v(n_45220_40040))
let min_45220_42840 = minimum(v(n_45220_42840))
let min_45220_45640 = minimum(v(n_45220_45640))
let min_45220_48440 = minimum(v(n_45220_48440))
let min_45220_51240 = minimum(v(n_45220_51240))
let min_45600_40040 = minimum(v(n_45600_40040))
let min_45600_42840 = minimum(v(n_45600_42840))
let min_45600_45640 = minimum(v(n_45600_45640))
let min_45600_48440 = minimum(v(n_45600_48440))
let min_45600_51240 = minimum(v(n_45600_51240))
let min_46360_40040 = minimum(v(n_46360_40040))
let min_46360_42840 = minimum(v(n_46360_42840))
let min_46360_45640 = minimum(v(n_46360_45640))
let min_46360_48440 = minimum(v(n_46360_48440))
let min_46360_51240 = minimum(v(n_46360_51240))
let min_46740_40040 = minimum(v(n_46740_40040))
let min_46740_42840 = minimum(v(n_46740_42840))
let min_46740_45640 = minimum(v(n_46740_45640))
let min_46740_48440 = minimum(v(n_46740_48440))
let min_46740_51240 = minimum(v(n_46740_51240))
let min_47120_40040 = minimum(v(n_47120_40040))
let min_47120_42840 = minimum(v(n_47120_42840))
let min_47120_45640 = minimum(v(n_47120_45640))
let min_47120_48440 = minimum(v(n_47120_48440))
let min_47120_51240 = minimum(v(n_47120_51240))
let min_47500_40040 = minimum(v(n_47500_40040))
let min_47500_42840 = minimum(v(n_47500_42840))
let min_47500_45640 = minimum(v(n_47500_45640))
let min_47500_48440 = minimum(v(n_47500_48440))
let min_47500_51240 = minimum(v(n_47500_51240))
let min_47880_40040 = minimum(v(n_47880_40040))
let min_47880_42840 = minimum(v(n_47880_42840))
let min_47880_45640 = minimum(v(n_47880_45640))
let min_47880_48440 = minimum(v(n_47880_48440))
let min_47880_51240 = minimum(v(n_47880_51240))
let min_48260_40040 = minimum(v(n_48260_40040))
let min_48260_42840 = minimum(v(n_48260_42840))
let min_48260_45640 = minimum(v(n_48260_45640))
let min_48260_48440 = minimum(v(n_48260_48440))
let min_48260_51240 = minimum(v(n_48260_51240))
let min_48640_40040 = minimum(v(n_48640_40040))
let min_48640_42840 = minimum(v(n_48640_42840))
let min_48640_45640 = minimum(v(n_48640_45640))
let min_48640_48440 = minimum(v(n_48640_48440))
let min_48640_51240 = minimum(v(n_48640_51240))
let min_49400_40040 = minimum(v(n_49400_40040))
let min_49400_42840 = minimum(v(n_49400_42840))
let min_49400_45640 = minimum(v(n_49400_45640))
let min_49400_48440 = minimum(v(n_49400_48440))
let min_49400_51240 = minimum(v(n_49400_51240))
let min_49780_40040 = minimum(v(n_49780_40040))
let min_49780_42840 = minimum(v(n_49780_42840))
let min_49780_45640 = minimum(v(n_49780_45640))
let min_49780_48440 = minimum(v(n_49780_48440))
let min_49780_51240 = minimum(v(n_49780_51240))
let min_50160_40040 = minimum(v(n_50160_40040))
let min_50160_42840 = minimum(v(n_50160_42840))
let min_50160_45640 = minimum(v(n_50160_45640))
let min_50160_48440 = minimum(v(n_50160_48440))
let min_50160_51240 = minimum(v(n_50160_51240))
let min_50540_40040 = minimum(v(n_50540_40040))
let min_50540_42840 = minimum(v(n_50540_42840))
let min_50540_45640 = minimum(v(n_50540_45640))
let min_50540_48440 = minimum(v(n_50540_48440))
let min_50540_51240 = minimum(v(n_50540_51240))
let min_51300_40040 = minimum(v(n_51300_40040))
let min_51300_42840 = minimum(v(n_51300_42840))
let min_51300_45640 = minimum(v(n_51300_45640))
let min_51300_48440 = minimum(v(n_51300_48440))
let min_51300_51240 = minimum(v(n_51300_51240))
let min_51680_40040 = minimum(v(n_51680_40040))
let min_51680_42840 = minimum(v(n_51680_42840))
let min_51680_45640 = minimum(v(n_51680_45640))
let min_51680_48440 = minimum(v(n_51680_48440))
let min_51680_51240 = minimum(v(n_51680_51240))
let min_52440_40040 = minimum(v(n_52440_40040))
let min_52440_42840 = minimum(v(n_52440_42840))
let min_52440_45640 = minimum(v(n_52440_45640))
let min_52440_48440 = minimum(v(n_52440_48440))
let min_52440_51240 = minimum(v(n_52440_51240))
let min_52820_40040 = minimum(v(n_52820_40040))
let min_52820_42840 = minimum(v(n_52820_42840))
let min_52820_45640 = minimum(v(n_52820_45640))
let min_52820_48440 = minimum(v(n_52820_48440))
let min_52820_51240 = minimum(v(n_52820_51240))
let min_53580_40040 = minimum(v(n_53580_40040))
let min_53580_42840 = minimum(v(n_53580_42840))
let min_53580_45640 = minimum(v(n_53580_45640))
let min_53580_48440 = minimum(v(n_53580_48440))
let min_53580_51240 = minimum(v(n_53580_51240))
let min_53960_40040 = minimum(v(n_53960_40040))
let min_53960_42840 = minimum(v(n_53960_42840))
let min_53960_45640 = minimum(v(n_53960_45640))
let min_53960_48440 = minimum(v(n_53960_48440))
let min_53960_51240 = minimum(v(n_53960_51240))
let min_54340_40040 = minimum(v(n_54340_40040))
let min_54340_42840 = minimum(v(n_54340_42840))
let min_54340_45640 = minimum(v(n_54340_45640))
let min_54340_48440 = minimum(v(n_54340_48440))
let min_54340_51240 = minimum(v(n_54340_51240))
let min_54720_40040 = minimum(v(n_54720_40040))
let min_54720_42840 = minimum(v(n_54720_42840))
let min_54720_45640 = minimum(v(n_54720_45640))
let min_54720_48440 = minimum(v(n_54720_48440))
let min_54720_51240 = minimum(v(n_54720_51240))
let min_55100_40040 = minimum(v(n_55100_40040))
let min_55100_42840 = minimum(v(n_55100_42840))
let min_55100_45640 = minimum(v(n_55100_45640))
let min_55100_48440 = minimum(v(n_55100_48440))
let min_55100_51240 = minimum(v(n_55100_51240))
* now write(append) all minimums to a file. ">>" means append:
print min_40660_40040 >> minimums
print min_40660_42840 >> minimums
print min_40660_45640 >> minimums
print min_40660_48440 >> minimums
print min_40660_51240 >> minimums
print min_41040_40040 >> minimums
print min_41040_42840 >> minimums
print min_41040_45640 >> minimums
print min_41040_48440 >> minimums
print min_41040_51240 >> minimums
print min_42180_40040 >> minimums
print min_42180_42840 >> minimums
print min_42180_45640 >> minimums
print min_42180_48440 >> minimums
print min_42180_51240 >> minimums
print min_42560_40040 >> minimums
print min_42560_42840 >> minimums
print min_42560_45640 >> minimums
print min_42560_48440 >> minimums
print min_42560_51240 >> minimums
print min_42940_40040 >> minimums
print min_42940_42840 >> minimums
print min_42940_45640 >> minimums
print min_42940_48440 >> minimums
print min_42940_51240 >> minimums
print min_43700_40040 >> minimums
print min_43700_42840 >> minimums
print min_43700_45640 >> minimums
print min_43700_48440 >> minimums
print min_43700_51240 >> minimums
print min_44080_40040 >> minimums
print min_44080_42840 >> minimums
print min_44080_45640 >> minimums
print min_44080_48440 >> minimums
print min_44080_51240 >> minimums
print min_44840_40040 >> minimums
print min_44840_42840 >> minimums
print min_44840_45640 >> minimums
print min_44840_48440 >> minimums
print min_44840_51240 >> minimums
print min_45220_40040 >> minimums
print min_45220_42840 >> minimums
print min_45220_45640 >> minimums
print min_45220_48440 >> minimums
print min_45220_51240 >> minimums
print min_45600_40040 >> minimums
print min_45600_42840 >> minimums
print min_45600_45640 >> minimums
print min_45600_48440 >> minimums
print min_45600_51240 >> minimums
print min_46360_40040 >> minimums
print min_46360_42840 >> minimums
print min_46360_45640 >> minimums
print min_46360_48440 >> minimums
print min_46360_51240 >> minimums
print min_46740_40040 >> minimums
print min_46740_42840 >> minimums
print min_46740_45640 >> minimums
print min_46740_48440 >> minimums
print min_46740_51240 >> minimums
print min_47120_40040 >> minimums
print min_47120_42840 >> minimums
print min_47120_45640 >> minimums
print min_47120_48440 >> minimums
print min_47120_51240 >> minimums
print min_47500_40040 >> minimums
print min_47500_42840 >> minimums
print min_47500_45640 >> minimums
print min_47500_48440 >> minimums
print min_47500_51240 >> minimums
print min_47880_40040 >> minimums
print min_47880_42840 >> minimums
print min_47880_45640 >> minimums
print min_47880_48440 >> minimums
print min_47880_51240 >> minimums
print min_48260_40040 >> minimums
print min_48260_42840 >> minimums
print min_48260_45640 >> minimums
print min_48260_48440 >> minimums
print min_48260_51240 >> minimums
print min_48640_40040 >> minimums
print min_48640_42840 >> minimums
print min_48640_45640 >> minimums
print min_48640_48440 >> minimums
print min_48640_51240 >> minimums
print min_49400_40040 >> minimums
print min_49400_42840 >> minimums
print min_49400_45640 >> minimums
print min_49400_48440 >> minimums
print min_49400_51240 >> minimums
print min_49780_40040 >> minimums
print min_49780_42840 >> minimums
print min_49780_45640 >> minimums
print min_49780_48440 >> minimums
print min_49780_51240 >> minimums
print min_50160_40040 >> minimums
print min_50160_42840 >> minimums
print min_50160_45640 >> minimums
print min_50160_48440 >> minimums
print min_50160_51240 >> minimums
print min_50540_40040 >> minimums
print min_50540_42840 >> minimums
print min_50540_45640 >> minimums
print min_50540_48440 >> minimums
print min_50540_51240 >> minimums
print min_51300_40040 >> minimums
print min_51300_42840 >> minimums
print min_51300_45640 >> minimums
print min_51300_48440 >> minimums
print min_51300_51240 >> minimums
print min_51680_40040 >> minimums
print min_51680_42840 >> minimums
print min_51680_45640 >> minimums
print min_51680_48440 >> minimums
print min_51680_51240 >> minimums
print min_52440_40040 >> minimums
print min_52440_42840 >> minimums
print min_52440_45640 >> minimums
print min_52440_48440 >> minimums
print min_52440_51240 >> minimums
print min_52820_40040 >> minimums
print min_52820_42840 >> minimums
print min_52820_45640 >> minimums
print min_52820_48440 >> minimums
print min_52820_51240 >> minimums
print min_53580_40040 >> minimums
print min_53580_42840 >> minimums
print min_53580_45640 >> minimums
print min_53580_48440 >> minimums
print min_53580_51240 >> minimums
print min_53960_40040 >> minimums
print min_53960_42840 >> minimums
print min_53960_45640 >> minimums
print min_53960_48440 >> minimums
print min_53960_51240 >> minimums
print min_54340_40040 >> minimums
print min_54340_42840 >> minimums
print min_54340_45640 >> minimums
print min_54340_48440 >> minimums
print min_54340_51240 >> minimums
print min_54720_40040 >> minimums
print min_54720_42840 >> minimums
print min_54720_45640 >> minimums
print min_54720_48440 >> minimums
print min_54720_51240 >> minimums
print min_55100_40040 >> minimums
print min_55100_42840 >> minimums
print min_55100_45640 >> minimums
print min_55100_48440 >> minimums
print min_55100_51240 >> minimums

exit
.endc