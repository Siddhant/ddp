.title 1-layer Power Grid for b02.points
* resistance segment model:
.subckt Rseg 1 3
R1 1 2 0.583
L1 2 3 0.003n
C1 1 0 0.25e-12
C2 3 0 0.25e-12
.ends
* the horizontal resistors:
X1 n_40280_40040 n_40660_40040 Rseg
X2 n_40660_40040 n_41420_40040 Rseg
X3 n_41420_40040 n_41800_40040 Rseg
X4 n_41800_40040 n_42180_40040 Rseg
X5 n_42180_40040 n_42560_40040 Rseg
X6 n_42560_40040 n_42940_40040 Rseg
X7 n_42940_40040 n_43700_40040 Rseg
X8 n_43700_40040 n_44080_40040 Rseg
X9 n_44080_40040 n_44460_40040 Rseg
X10 n_44460_40040 n_44840_40040 Rseg
X11 n_44840_40040 n_45220_40040 Rseg
X12 n_45220_40040 n_45600_40040 Rseg
X13 n_45600_40040 n_45980_40040 Rseg
X14 n_45980_40040 n_46740_40040 Rseg
X15 n_46740_40040 n_47120_40040 Rseg
X16 n_47120_40040 n_47500_40040 Rseg
X17 n_47500_40040 n_48260_40040 Rseg
X18 n_48260_40040 n_48640_40040 Rseg
X19 n_48640_40040 n_49020_40040 Rseg
X20 n_49020_40040 n_49400_40040 Rseg
X21 n_49400_40040 n_50540_40040 Rseg
X22 n_50540_40040 n_50920_40040 Rseg
X23 n_50920_40040 n_51300_40040 Rseg
X24 n_51300_40040 n_51680_40040 Rseg
X25 n_51680_40040 n_53200_40040 Rseg
X26 n_40280_42840 n_40660_42840 Rseg
X27 n_40660_42840 n_41420_42840 Rseg
X28 n_41420_42840 n_41800_42840 Rseg
X29 n_41800_42840 n_42180_42840 Rseg
X30 n_42180_42840 n_42560_42840 Rseg
X31 n_42560_42840 n_42940_42840 Rseg
X32 n_42940_42840 n_43700_42840 Rseg
X33 n_43700_42840 n_44080_42840 Rseg
X34 n_44080_42840 n_44460_42840 Rseg
X35 n_44460_42840 n_44840_42840 Rseg
X36 n_44840_42840 n_45220_42840 Rseg
X37 n_45220_42840 n_45600_42840 Rseg
X38 n_45600_42840 n_45980_42840 Rseg
X39 n_45980_42840 n_46740_42840 Rseg
X40 n_46740_42840 n_47120_42840 Rseg
X41 n_47120_42840 n_47500_42840 Rseg
X42 n_47500_42840 n_48260_42840 Rseg
X43 n_48260_42840 n_48640_42840 Rseg
X44 n_48640_42840 n_49020_42840 Rseg
X45 n_49020_42840 n_49400_42840 Rseg
X46 n_49400_42840 n_50540_42840 Rseg
X47 n_50540_42840 n_50920_42840 Rseg
X48 n_50920_42840 n_51300_42840 Rseg
X49 n_51300_42840 n_51680_42840 Rseg
X50 n_51680_42840 n_53200_42840 Rseg
X51 n_40280_45640 n_40660_45640 Rseg
X52 n_40660_45640 n_41420_45640 Rseg
X53 n_41420_45640 n_41800_45640 Rseg
X54 n_41800_45640 n_42180_45640 Rseg
X55 n_42180_45640 n_42560_45640 Rseg
X56 n_42560_45640 n_42940_45640 Rseg
X57 n_42940_45640 n_43700_45640 Rseg
X58 n_43700_45640 n_44080_45640 Rseg
X59 n_44080_45640 n_44460_45640 Rseg
X60 n_44460_45640 n_44840_45640 Rseg
X61 n_44840_45640 n_45220_45640 Rseg
X62 n_45220_45640 n_45600_45640 Rseg
X63 n_45600_45640 n_45980_45640 Rseg
X64 n_45980_45640 n_46740_45640 Rseg
X65 n_46740_45640 n_47120_45640 Rseg
X66 n_47120_45640 n_47500_45640 Rseg
X67 n_47500_45640 n_48260_45640 Rseg
X68 n_48260_45640 n_48640_45640 Rseg
X69 n_48640_45640 n_49020_45640 Rseg
X70 n_49020_45640 n_49400_45640 Rseg
X71 n_49400_45640 n_50540_45640 Rseg
X72 n_50540_45640 n_50920_45640 Rseg
X73 n_50920_45640 n_51300_45640 Rseg
X74 n_51300_45640 n_51680_45640 Rseg
X75 n_51680_45640 n_53200_45640 Rseg
* the vertical resistors:
X76 n_40280_40040 n_40280_42840 Rseg
X77 n_40280_42840 n_40280_45640 Rseg
X78 n_40660_40040 n_40660_42840 Rseg
X79 n_40660_42840 n_40660_45640 Rseg
X80 n_41420_40040 n_41420_42840 Rseg
X81 n_41420_42840 n_41420_45640 Rseg
X82 n_41800_40040 n_41800_42840 Rseg
X83 n_41800_42840 n_41800_45640 Rseg
X84 n_42180_40040 n_42180_42840 Rseg
X85 n_42180_42840 n_42180_45640 Rseg
X86 n_42560_40040 n_42560_42840 Rseg
X87 n_42560_42840 n_42560_45640 Rseg
X88 n_42940_40040 n_42940_42840 Rseg
X89 n_42940_42840 n_42940_45640 Rseg
X90 n_43700_40040 n_43700_42840 Rseg
X91 n_43700_42840 n_43700_45640 Rseg
X92 n_44080_40040 n_44080_42840 Rseg
X93 n_44080_42840 n_44080_45640 Rseg
X94 n_44460_40040 n_44460_42840 Rseg
X95 n_44460_42840 n_44460_45640 Rseg
X96 n_44840_40040 n_44840_42840 Rseg
X97 n_44840_42840 n_44840_45640 Rseg
X98 n_45220_40040 n_45220_42840 Rseg
X99 n_45220_42840 n_45220_45640 Rseg
X100 n_45600_40040 n_45600_42840 Rseg
X101 n_45600_42840 n_45600_45640 Rseg
X102 n_45980_40040 n_45980_42840 Rseg
X103 n_45980_42840 n_45980_45640 Rseg
X104 n_46740_40040 n_46740_42840 Rseg
X105 n_46740_42840 n_46740_45640 Rseg
X106 n_47120_40040 n_47120_42840 Rseg
X107 n_47120_42840 n_47120_45640 Rseg
X108 n_47500_40040 n_47500_42840 Rseg
X109 n_47500_42840 n_47500_45640 Rseg
X110 n_48260_40040 n_48260_42840 Rseg
X111 n_48260_42840 n_48260_45640 Rseg
X112 n_48640_40040 n_48640_42840 Rseg
X113 n_48640_42840 n_48640_45640 Rseg
X114 n_49020_40040 n_49020_42840 Rseg
X115 n_49020_42840 n_49020_45640 Rseg
X116 n_49400_40040 n_49400_42840 Rseg
X117 n_49400_42840 n_49400_45640 Rseg
X118 n_50540_40040 n_50540_42840 Rseg
X119 n_50540_42840 n_50540_45640 Rseg
X120 n_50920_40040 n_50920_42840 Rseg
X121 n_50920_42840 n_50920_45640 Rseg
X122 n_51300_40040 n_51300_42840 Rseg
X123 n_51300_42840 n_51300_45640 Rseg
X124 n_51680_40040 n_51680_42840 Rseg
X125 n_51680_42840 n_51680_45640 Rseg
X126 n_53200_40040 n_53200_42840 Rseg
X127 n_53200_42840 n_53200_45640 Rseg
* voltage source is placed at (x_min, y_min)
Vin n_40280_40040 0 DC 1.0

I1 n_51300_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I2 n_53200_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I3 n_51680_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I4 n_41420_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I5 n_42560_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I6 n_42940_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I7 n_44080_45640 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I8 n_49020_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I9 n_47120_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I10 n_44840_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I11 n_47500_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I12 n_50540_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I13 n_49400_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I14 n_48640_42840 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I15 n_44460_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I16 n_42940_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I17 n_42180_40040 0 PWL(0ps 0uA 30ps 0uA 31ps 30uA 59ps 30uA 60ps 0uA)
I18 n_51300_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I19 n_44080_45640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I20 n_49020_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I21 n_47120_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I22 n_47500_42840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I23 n_48640_42840 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I24 n_44460_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I25 n_42940_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I26 n_42180_40040 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I27 n_49400_45640 0 PWL(2000ps 0uA 2030ps 0uA 2031ps 30uA 2059ps 30uA 2060ps 0uA)
I28 n_51300_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I29 n_53200_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I30 n_41420_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I31 n_42560_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I32 n_45980_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I33 n_45220_45640 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I34 n_49020_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I35 n_47120_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I36 n_43700_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I37 n_48640_42840 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I38 n_44460_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I39 n_40660_40040 0 PWL(4000ps 0uA 4030ps 0uA 4031ps 30uA 4059ps 30uA 4060ps 0uA)
I40 n_51680_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I41 n_45980_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I42 n_42940_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I43 n_43700_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I44 n_44840_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I45 n_50540_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I46 n_49400_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I47 n_46740_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I48 n_48640_42840 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I49 n_44460_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I50 n_40660_40040 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I51 n_49400_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I52 n_48260_45640 0 PWL(6000ps 0uA 6030ps 0uA 6031ps 30uA 6059ps 30uA 6060ps 0uA)
I53 n_51300_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I54 n_51680_42840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I55 n_40660_45640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I56 n_41800_45640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I57 n_45980_45640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I58 n_45220_45640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I59 n_49020_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I60 n_45600_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I61 n_44840_42840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I62 n_47500_42840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I63 n_50540_42840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I64 n_49400_42840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I65 n_46740_45640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I66 n_48640_42840 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I67 n_44460_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I68 n_42940_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I69 n_42180_40040 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I70 n_48260_45640 0 PWL(8000ps 0uA 8030ps 0uA 8031ps 30uA 8059ps 30uA 8060ps 0uA)
I71 n_51300_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I72 n_53200_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I73 n_51680_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I74 n_41420_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I75 n_40280_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I76 n_45220_45640 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I77 n_49020_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I78 n_45600_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I79 n_43700_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I80 n_50540_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I81 n_49400_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I82 n_48640_42840 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I83 n_44460_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I84 n_42940_40040 0 PWL(10000ps 0uA 10030ps 0uA 10031ps 30uA 10059ps 30uA 10060ps 0uA)
I85 n_51300_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I86 n_51680_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I87 n_49020_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I88 n_45600_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I89 n_43700_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I90 n_44840_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I91 n_47500_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I92 n_50540_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I93 n_49400_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I94 n_48640_42840 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I95 n_44460_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I96 n_40660_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I97 n_42180_40040 0 PWL(12000ps 0uA 12030ps 0uA 12031ps 30uA 12059ps 30uA 12060ps 0uA)
I98 n_42560_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I99 n_40280_42840 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I100 n_40660_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I101 n_41800_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I102 n_45980_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I103 n_42940_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I104 n_45220_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I105 n_44080_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I106 n_47120_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I107 n_45600_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I108 n_42940_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I109 n_40660_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I110 n_42180_40040 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I111 n_49400_45640 0 PWL(14000ps 0uA 14030ps 0uA 14031ps 30uA 14059ps 30uA 14060ps 0uA)
I112 n_53200_40040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I113 n_51300_40040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I114 n_53200_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I115 n_51680_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I116 n_50920_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I117 n_53200_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I118 n_41420_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I119 n_42560_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I120 n_45220_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I121 n_44080_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I122 n_49020_40040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I123 n_47120_40040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I124 n_43700_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I125 n_44840_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I126 n_50540_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I127 n_46740_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I128 n_48640_42840 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I129 n_44460_40040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I130 n_42940_40040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I131 n_42180_40040 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
I132 n_48260_45640 0 PWL(16000ps 0uA 16030ps 0uA 16031ps 30uA 16059ps 30uA 16060ps 0uA)
.tran 1ps 20000ps
.control
run
* calculate minimum value of voltage at each node:
let min_40280_40040 = minimum(v(n_40280_40040))
let min_40280_42840 = minimum(v(n_40280_42840))
let min_40280_45640 = minimum(v(n_40280_45640))
let min_40660_40040 = minimum(v(n_40660_40040))
let min_40660_42840 = minimum(v(n_40660_42840))
let min_40660_45640 = minimum(v(n_40660_45640))
let min_41420_40040 = minimum(v(n_41420_40040))
let min_41420_42840 = minimum(v(n_41420_42840))
let min_41420_45640 = minimum(v(n_41420_45640))
let min_41800_40040 = minimum(v(n_41800_40040))
let min_41800_42840 = minimum(v(n_41800_42840))
let min_41800_45640 = minimum(v(n_41800_45640))
let min_42180_40040 = minimum(v(n_42180_40040))
let min_42180_42840 = minimum(v(n_42180_42840))
let min_42180_45640 = minimum(v(n_42180_45640))
let min_42560_40040 = minimum(v(n_42560_40040))
let min_42560_42840 = minimum(v(n_42560_42840))
let min_42560_45640 = minimum(v(n_42560_45640))
let min_42940_40040 = minimum(v(n_42940_40040))
let min_42940_42840 = minimum(v(n_42940_42840))
let min_42940_45640 = minimum(v(n_42940_45640))
let min_43700_40040 = minimum(v(n_43700_40040))
let min_43700_42840 = minimum(v(n_43700_42840))
let min_43700_45640 = minimum(v(n_43700_45640))
let min_44080_40040 = minimum(v(n_44080_40040))
let min_44080_42840 = minimum(v(n_44080_42840))
let min_44080_45640 = minimum(v(n_44080_45640))
let min_44460_40040 = minimum(v(n_44460_40040))
let min_44460_42840 = minimum(v(n_44460_42840))
let min_44460_45640 = minimum(v(n_44460_45640))
let min_44840_40040 = minimum(v(n_44840_40040))
let min_44840_42840 = minimum(v(n_44840_42840))
let min_44840_45640 = minimum(v(n_44840_45640))
let min_45220_40040 = minimum(v(n_45220_40040))
let min_45220_42840 = minimum(v(n_45220_42840))
let min_45220_45640 = minimum(v(n_45220_45640))
let min_45600_40040 = minimum(v(n_45600_40040))
let min_45600_42840 = minimum(v(n_45600_42840))
let min_45600_45640 = minimum(v(n_45600_45640))
let min_45980_40040 = minimum(v(n_45980_40040))
let min_45980_42840 = minimum(v(n_45980_42840))
let min_45980_45640 = minimum(v(n_45980_45640))
let min_46740_40040 = minimum(v(n_46740_40040))
let min_46740_42840 = minimum(v(n_46740_42840))
let min_46740_45640 = minimum(v(n_46740_45640))
let min_47120_40040 = minimum(v(n_47120_40040))
let min_47120_42840 = minimum(v(n_47120_42840))
let min_47120_45640 = minimum(v(n_47120_45640))
let min_47500_40040 = minimum(v(n_47500_40040))
let min_47500_42840 = minimum(v(n_47500_42840))
let min_47500_45640 = minimum(v(n_47500_45640))
let min_48260_40040 = minimum(v(n_48260_40040))
let min_48260_42840 = minimum(v(n_48260_42840))
let min_48260_45640 = minimum(v(n_48260_45640))
let min_48640_40040 = minimum(v(n_48640_40040))
let min_48640_42840 = minimum(v(n_48640_42840))
let min_48640_45640 = minimum(v(n_48640_45640))
let min_49020_40040 = minimum(v(n_49020_40040))
let min_49020_42840 = minimum(v(n_49020_42840))
let min_49020_45640 = minimum(v(n_49020_45640))
let min_49400_40040 = minimum(v(n_49400_40040))
let min_49400_42840 = minimum(v(n_49400_42840))
let min_49400_45640 = minimum(v(n_49400_45640))
let min_50540_40040 = minimum(v(n_50540_40040))
let min_50540_42840 = minimum(v(n_50540_42840))
let min_50540_45640 = minimum(v(n_50540_45640))
let min_50920_40040 = minimum(v(n_50920_40040))
let min_50920_42840 = minimum(v(n_50920_42840))
let min_50920_45640 = minimum(v(n_50920_45640))
let min_51300_40040 = minimum(v(n_51300_40040))
let min_51300_42840 = minimum(v(n_51300_42840))
let min_51300_45640 = minimum(v(n_51300_45640))
let min_51680_40040 = minimum(v(n_51680_40040))
let min_51680_42840 = minimum(v(n_51680_42840))
let min_51680_45640 = minimum(v(n_51680_45640))
let min_53200_40040 = minimum(v(n_53200_40040))
let min_53200_42840 = minimum(v(n_53200_42840))
let min_53200_45640 = minimum(v(n_53200_45640))
* now write(append) all minimums to a file. ">>" means append:
print min_40280_40040 >> minimums
print min_40280_42840 >> minimums
print min_40280_45640 >> minimums
print min_40660_40040 >> minimums
print min_40660_42840 >> minimums
print min_40660_45640 >> minimums
print min_41420_40040 >> minimums
print min_41420_42840 >> minimums
print min_41420_45640 >> minimums
print min_41800_40040 >> minimums
print min_41800_42840 >> minimums
print min_41800_45640 >> minimums
print min_42180_40040 >> minimums
print min_42180_42840 >> minimums
print min_42180_45640 >> minimums
print min_42560_40040 >> minimums
print min_42560_42840 >> minimums
print min_42560_45640 >> minimums
print min_42940_40040 >> minimums
print min_42940_42840 >> minimums
print min_42940_45640 >> minimums
print min_43700_40040 >> minimums
print min_43700_42840 >> minimums
print min_43700_45640 >> minimums
print min_44080_40040 >> minimums
print min_44080_42840 >> minimums
print min_44080_45640 >> minimums
print min_44460_40040 >> minimums
print min_44460_42840 >> minimums
print min_44460_45640 >> minimums
print min_44840_40040 >> minimums
print min_44840_42840 >> minimums
print min_44840_45640 >> minimums
print min_45220_40040 >> minimums
print min_45220_42840 >> minimums
print min_45220_45640 >> minimums
print min_45600_40040 >> minimums
print min_45600_42840 >> minimums
print min_45600_45640 >> minimums
print min_45980_40040 >> minimums
print min_45980_42840 >> minimums
print min_45980_45640 >> minimums
print min_46740_40040 >> minimums
print min_46740_42840 >> minimums
print min_46740_45640 >> minimums
print min_47120_40040 >> minimums
print min_47120_42840 >> minimums
print min_47120_45640 >> minimums
print min_47500_40040 >> minimums
print min_47500_42840 >> minimums
print min_47500_45640 >> minimums
print min_48260_40040 >> minimums
print min_48260_42840 >> minimums
print min_48260_45640 >> minimums
print min_48640_40040 >> minimums
print min_48640_42840 >> minimums
print min_48640_45640 >> minimums
print min_49020_40040 >> minimums
print min_49020_42840 >> minimums
print min_49020_45640 >> minimums
print min_49400_40040 >> minimums
print min_49400_42840 >> minimums
print min_49400_45640 >> minimums
print min_50540_40040 >> minimums
print min_50540_42840 >> minimums
print min_50540_45640 >> minimums
print min_50920_40040 >> minimums
print min_50920_42840 >> minimums
print min_50920_45640 >> minimums
print min_51300_40040 >> minimums
print min_51300_42840 >> minimums
print min_51300_45640 >> minimums
print min_51680_40040 >> minimums
print min_51680_42840 >> minimums
print min_51680_45640 >> minimums
print min_53200_40040 >> minimums
print min_53200_42840 >> minimums
print min_53200_45640 >> minimums

exit
.endc